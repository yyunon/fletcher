-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Interconnect_pkg.all;

entity Abs_kernel_Mantle is
  generic (
    INDEX_WIDTH        : integer := 32;
    TAG_WIDTH          : integer := 1;
    BUS_ADDR_WIDTH     : integer := 64;
    BUS_DATA_WIDTH     : integer := 512;
    BUS_LEN_WIDTH      : integer := 8;
    BUS_BURST_STEP_LEN : integer := 1;
    BUS_BURST_MAX_LEN  : integer := 16
  );
  port (
    bcd_clk            : in  std_logic;
    bcd_reset          : in  std_logic;
    kcd_clk            : in  std_logic;
    kcd_reset          : in  std_logic;
    mmio_awvalid       : in  std_logic;
    mmio_awready       : out std_logic;
    mmio_awaddr        : in  std_logic_vector(31 downto 0);
    mmio_wvalid        : in  std_logic;
    mmio_wready        : out std_logic;
    mmio_wdata         : in  std_logic_vector(31 downto 0);
    mmio_wstrb         : in  std_logic_vector(3 downto 0);
    mmio_bvalid        : out std_logic;
    mmio_bready        : in  std_logic;
    mmio_bresp         : out std_logic_vector(1 downto 0);
    mmio_arvalid       : in  std_logic;
    mmio_arready       : out std_logic;
    mmio_araddr        : in  std_logic_vector(31 downto 0);
    mmio_rvalid        : out std_logic;
    mmio_rready        : in  std_logic;
    mmio_rdata         : out std_logic_vector(31 downto 0);
    mmio_rresp         : out std_logic_vector(1 downto 0);
    rd_mst_rreq_valid  : out std_logic;
    rd_mst_rreq_ready  : in  std_logic;
    rd_mst_rreq_addr   : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    rd_mst_rreq_len    : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    rd_mst_rdat_valid  : in  std_logic;
    rd_mst_rdat_ready  : out std_logic;
    rd_mst_rdat_data   : in  std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    rd_mst_rdat_last   : in  std_logic;
    wr_mst_wreq_valid  : out std_logic;
    wr_mst_wreq_ready  : in  std_logic;
    wr_mst_wreq_addr   : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    wr_mst_wreq_len    : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    wr_mst_wdat_valid  : out std_logic;
    wr_mst_wdat_ready  : in  std_logic;
    wr_mst_wdat_data   : out std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    wr_mst_wdat_strobe : out std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
    wr_mst_wdat_last   : out std_logic
  );
end entity;

architecture Implementation of Abs_kernel_Mantle is
  component Abs_kernel_Nucleus is
    generic (
      INDEX_WIDTH                     : integer := 32;
      TAG_WIDTH                       : integer := 1;
      BATCHIN_VECTORS_BUS_ADDR_WIDTH  : integer := 64;
      BATCHOUT_VECTORS_BUS_ADDR_WIDTH : integer := 64
    );
    port (
      kcd_clk                       : in  std_logic;
      kcd_reset                     : in  std_logic;
      mmio_awvalid                  : in  std_logic;
      mmio_awready                  : out std_logic;
      mmio_awaddr                   : in  std_logic_vector(31 downto 0);
      mmio_wvalid                   : in  std_logic;
      mmio_wready                   : out std_logic;
      mmio_wdata                    : in  std_logic_vector(31 downto 0);
      mmio_wstrb                    : in  std_logic_vector(3 downto 0);
      mmio_bvalid                   : out std_logic;
      mmio_bready                   : in  std_logic;
      mmio_bresp                    : out std_logic_vector(1 downto 0);
      mmio_arvalid                  : in  std_logic;
      mmio_arready                  : out std_logic;
      mmio_araddr                   : in  std_logic_vector(31 downto 0);
      mmio_rvalid                   : out std_logic;
      mmio_rready                   : in  std_logic;
      mmio_rdata                    : out std_logic_vector(31 downto 0);
      mmio_rresp                    : out std_logic_vector(1 downto 0);
      BatchIn_vectors_valid         : in  std_logic;
      BatchIn_vectors_ready         : out std_logic;
      BatchIn_vectors_dvalid        : in  std_logic;
      BatchIn_vectors_last          : in  std_logic;
      BatchIn_vectors               : in  std_logic_vector(63 downto 0);
      BatchIn_vectors_unl_valid     : in  std_logic;
      BatchIn_vectors_unl_ready     : out std_logic;
      BatchIn_vectors_unl_tag       : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      BatchIn_vectors_cmd_valid     : out std_logic;
      BatchIn_vectors_cmd_ready     : in  std_logic;
      BatchIn_vectors_cmd_firstIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      BatchIn_vectors_cmd_lastIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      BatchIn_vectors_cmd_ctrl      : out std_logic_vector(BATCHIN_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
      BatchIn_vectors_cmd_tag       : out std_logic_vector(TAG_WIDTH-1 downto 0);
      BatchOut_vectors_valid        : out std_logic;
      BatchOut_vectors_ready        : in  std_logic;
      BatchOut_vectors_dvalid       : out std_logic;
      BatchOut_vectors_last         : out std_logic;
      BatchOut_vectors              : out std_logic_vector(63 downto 0);
      BatchOut_vectors_unl_valid    : in  std_logic;
      BatchOut_vectors_unl_ready    : out std_logic;
      BatchOut_vectors_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      BatchOut_vectors_cmd_valid    : out std_logic;
      BatchOut_vectors_cmd_ready    : in  std_logic;
      BatchOut_vectors_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      BatchOut_vectors_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      BatchOut_vectors_cmd_ctrl     : out std_logic_vector(BATCHOUT_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
      BatchOut_vectors_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Abs_kernel_BatchIn is
    generic (
      INDEX_WIDTH                        : integer := 32;
      TAG_WIDTH                          : integer := 1;
      BATCHIN_VECTORS_BUS_ADDR_WIDTH     : integer := 64;
      BATCHIN_VECTORS_BUS_DATA_WIDTH     : integer := 512;
      BATCHIN_VECTORS_BUS_LEN_WIDTH      : integer := 8;
      BATCHIN_VECTORS_BUS_BURST_STEP_LEN : integer := 1;
      BATCHIN_VECTORS_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                        : in  std_logic;
      bcd_reset                      : in  std_logic;
      kcd_clk                        : in  std_logic;
      kcd_reset                      : in  std_logic;
      BatchIn_vectors_valid          : out std_logic;
      BatchIn_vectors_ready          : in  std_logic;
      BatchIn_vectors_dvalid         : out std_logic;
      BatchIn_vectors_last           : out std_logic;
      BatchIn_vectors                : out std_logic_vector(63 downto 0);
      BatchIn_vectors_bus_rreq_valid : out std_logic;
      BatchIn_vectors_bus_rreq_ready : in  std_logic;
      BatchIn_vectors_bus_rreq_addr  : out std_logic_vector(BATCHIN_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
      BatchIn_vectors_bus_rreq_len   : out std_logic_vector(BATCHIN_VECTORS_BUS_LEN_WIDTH-1 downto 0);
      BatchIn_vectors_bus_rdat_valid : in  std_logic;
      BatchIn_vectors_bus_rdat_ready : out std_logic;
      BatchIn_vectors_bus_rdat_data  : in  std_logic_vector(BATCHIN_VECTORS_BUS_DATA_WIDTH-1 downto 0);
      BatchIn_vectors_bus_rdat_last  : in  std_logic;
      BatchIn_vectors_cmd_valid      : in  std_logic;
      BatchIn_vectors_cmd_ready      : out std_logic;
      BatchIn_vectors_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      BatchIn_vectors_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      BatchIn_vectors_cmd_ctrl       : in  std_logic_vector(BATCHIN_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
      BatchIn_vectors_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      BatchIn_vectors_unl_valid      : out std_logic;
      BatchIn_vectors_unl_ready      : in  std_logic;
      BatchIn_vectors_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Abs_kernel_BatchOut is
    generic (
      INDEX_WIDTH                         : integer := 32;
      TAG_WIDTH                           : integer := 1;
      BATCHOUT_VECTORS_BUS_ADDR_WIDTH     : integer := 64;
      BATCHOUT_VECTORS_BUS_DATA_WIDTH     : integer := 512;
      BATCHOUT_VECTORS_BUS_LEN_WIDTH      : integer := 8;
      BATCHOUT_VECTORS_BUS_BURST_STEP_LEN : integer := 1;
      BATCHOUT_VECTORS_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                          : in  std_logic;
      bcd_reset                        : in  std_logic;
      kcd_clk                          : in  std_logic;
      kcd_reset                        : in  std_logic;
      BatchOut_vectors_valid           : in  std_logic;
      BatchOut_vectors_ready           : out std_logic;
      BatchOut_vectors_dvalid          : in  std_logic;
      BatchOut_vectors_last            : in  std_logic;
      BatchOut_vectors                 : in  std_logic_vector(63 downto 0);
      BatchOut_vectors_bus_wreq_valid  : out std_logic;
      BatchOut_vectors_bus_wreq_ready  : in  std_logic;
      BatchOut_vectors_bus_wreq_addr   : out std_logic_vector(BATCHOUT_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
      BatchOut_vectors_bus_wreq_len    : out std_logic_vector(BATCHOUT_VECTORS_BUS_LEN_WIDTH-1 downto 0);
      BatchOut_vectors_bus_wdat_valid  : out std_logic;
      BatchOut_vectors_bus_wdat_ready  : in  std_logic;
      BatchOut_vectors_bus_wdat_data   : out std_logic_vector(BATCHOUT_VECTORS_BUS_DATA_WIDTH-1 downto 0);
      BatchOut_vectors_bus_wdat_strobe : out std_logic_vector(BATCHOUT_VECTORS_BUS_DATA_WIDTH/8-1 downto 0);
      BatchOut_vectors_bus_wdat_last   : out std_logic;
      BatchOut_vectors_cmd_valid       : in  std_logic;
      BatchOut_vectors_cmd_ready       : out std_logic;
      BatchOut_vectors_cmd_firstIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      BatchOut_vectors_cmd_lastIdx     : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      BatchOut_vectors_cmd_ctrl        : in  std_logic_vector(BATCHOUT_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
      BatchOut_vectors_cmd_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      BatchOut_vectors_unl_valid       : out std_logic;
      BatchOut_vectors_unl_ready       : in  std_logic;
      BatchOut_vectors_unl_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  signal Abs_kernel_Nucleus_inst_kcd_clk                           : std_logic;
  signal Abs_kernel_Nucleus_inst_kcd_reset                         : std_logic;

  signal Abs_kernel_Nucleus_inst_mmio_awvalid                      : std_logic;
  signal Abs_kernel_Nucleus_inst_mmio_awready                      : std_logic;
  signal Abs_kernel_Nucleus_inst_mmio_awaddr                       : std_logic_vector(31 downto 0);
  signal Abs_kernel_Nucleus_inst_mmio_wvalid                       : std_logic;
  signal Abs_kernel_Nucleus_inst_mmio_wready                       : std_logic;
  signal Abs_kernel_Nucleus_inst_mmio_wdata                        : std_logic_vector(31 downto 0);
  signal Abs_kernel_Nucleus_inst_mmio_wstrb                        : std_logic_vector(3 downto 0);
  signal Abs_kernel_Nucleus_inst_mmio_bvalid                       : std_logic;
  signal Abs_kernel_Nucleus_inst_mmio_bready                       : std_logic;
  signal Abs_kernel_Nucleus_inst_mmio_bresp                        : std_logic_vector(1 downto 0);
  signal Abs_kernel_Nucleus_inst_mmio_arvalid                      : std_logic;
  signal Abs_kernel_Nucleus_inst_mmio_arready                      : std_logic;
  signal Abs_kernel_Nucleus_inst_mmio_araddr                       : std_logic_vector(31 downto 0);
  signal Abs_kernel_Nucleus_inst_mmio_rvalid                       : std_logic;
  signal Abs_kernel_Nucleus_inst_mmio_rready                       : std_logic;
  signal Abs_kernel_Nucleus_inst_mmio_rdata                        : std_logic_vector(31 downto 0);
  signal Abs_kernel_Nucleus_inst_mmio_rresp                        : std_logic_vector(1 downto 0);

  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_valid             : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_ready             : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_dvalid            : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_last              : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchIn_vectors                   : std_logic_vector(63 downto 0);

  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_unl_valid         : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_unl_ready         : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_valid         : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_ready         : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_valid            : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_ready            : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_dvalid           : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_last             : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchOut_vectors                  : std_logic_vector(63 downto 0);

  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_unl_valid        : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_unl_ready        : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_unl_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_valid        : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_ready        : std_logic;
  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_ctrl         : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Abs_kernel_BatchIn_inst_bcd_clk                           : std_logic;
  signal Abs_kernel_BatchIn_inst_bcd_reset                         : std_logic;

  signal Abs_kernel_BatchIn_inst_kcd_clk                           : std_logic;
  signal Abs_kernel_BatchIn_inst_kcd_reset                         : std_logic;

  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_valid             : std_logic;
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_ready             : std_logic;
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_dvalid            : std_logic;
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_last              : std_logic;
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors                   : std_logic_vector(63 downto 0);

  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rreq_valid    : std_logic;
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rreq_ready    : std_logic;
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rreq_addr     : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rreq_len      : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rdat_valid    : std_logic;
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rdat_ready    : std_logic;
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rdat_data     : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rdat_last     : std_logic;

  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_valid         : std_logic;
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_ready         : std_logic;
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_unl_valid         : std_logic;
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_unl_ready         : std_logic;
  signal Abs_kernel_BatchIn_inst_BatchIn_vectors_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Abs_kernel_BatchOut_inst_bcd_clk                          : std_logic;
  signal Abs_kernel_BatchOut_inst_bcd_reset                        : std_logic;

  signal Abs_kernel_BatchOut_inst_kcd_clk                          : std_logic;
  signal Abs_kernel_BatchOut_inst_kcd_reset                        : std_logic;

  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_valid           : std_logic;
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_ready           : std_logic;
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_dvalid          : std_logic;
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_last            : std_logic;
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors                 : std_logic_vector(63 downto 0);

  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wreq_valid  : std_logic;
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wreq_ready  : std_logic;
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wreq_addr   : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wreq_len    : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_valid  : std_logic;
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_ready  : std_logic;
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_data   : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_strobe : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_last   : std_logic;

  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_valid       : std_logic;
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_ready       : std_logic;
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_ctrl        : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_unl_valid       : std_logic;
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_unl_ready       : std_logic;
  signal Abs_kernel_BatchOut_inst_BatchOut_vectors_unl_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal RDAW64DW512LW8BS1BM16_inst_bcd_clk                        : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_bcd_reset                      : std_logic;

  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid                 : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready                 : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr                  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_len                   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid                 : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready                 : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_data                  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_last                  : std_logic;

  signal WRAW64DW512LW8BS1BM16_inst_bcd_clk                        : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_bcd_reset                      : std_logic;

  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid                 : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready                 : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr                  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_len                   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid                 : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready                 : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_data                  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe                : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_last                  : std_logic;

  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid  : std_logic_vector(0 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready  : std_logic_vector(0 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr   : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len    : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid  : std_logic_vector(0 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready  : std_logic_vector(0 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data   : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last   : std_logic_vector(0 downto 0);

  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid  : std_logic_vector(0 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready  : std_logic_vector(0 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr   : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len    : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid  : std_logic_vector(0 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready  : std_logic_vector(0 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data   : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last   : std_logic_vector(0 downto 0);

begin
  Abs_kernel_Nucleus_inst : Abs_kernel_Nucleus
    generic map (
      INDEX_WIDTH                     => INDEX_WIDTH,
      TAG_WIDTH                       => TAG_WIDTH,
      BATCHIN_VECTORS_BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
      BATCHOUT_VECTORS_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH
    )
    port map (
      kcd_clk                       => Abs_kernel_Nucleus_inst_kcd_clk,
      kcd_reset                     => Abs_kernel_Nucleus_inst_kcd_reset,
      mmio_awvalid                  => Abs_kernel_Nucleus_inst_mmio_awvalid,
      mmio_awready                  => Abs_kernel_Nucleus_inst_mmio_awready,
      mmio_awaddr                   => Abs_kernel_Nucleus_inst_mmio_awaddr,
      mmio_wvalid                   => Abs_kernel_Nucleus_inst_mmio_wvalid,
      mmio_wready                   => Abs_kernel_Nucleus_inst_mmio_wready,
      mmio_wdata                    => Abs_kernel_Nucleus_inst_mmio_wdata,
      mmio_wstrb                    => Abs_kernel_Nucleus_inst_mmio_wstrb,
      mmio_bvalid                   => Abs_kernel_Nucleus_inst_mmio_bvalid,
      mmio_bready                   => Abs_kernel_Nucleus_inst_mmio_bready,
      mmio_bresp                    => Abs_kernel_Nucleus_inst_mmio_bresp,
      mmio_arvalid                  => Abs_kernel_Nucleus_inst_mmio_arvalid,
      mmio_arready                  => Abs_kernel_Nucleus_inst_mmio_arready,
      mmio_araddr                   => Abs_kernel_Nucleus_inst_mmio_araddr,
      mmio_rvalid                   => Abs_kernel_Nucleus_inst_mmio_rvalid,
      mmio_rready                   => Abs_kernel_Nucleus_inst_mmio_rready,
      mmio_rdata                    => Abs_kernel_Nucleus_inst_mmio_rdata,
      mmio_rresp                    => Abs_kernel_Nucleus_inst_mmio_rresp,
      BatchIn_vectors_valid         => Abs_kernel_Nucleus_inst_BatchIn_vectors_valid,
      BatchIn_vectors_ready         => Abs_kernel_Nucleus_inst_BatchIn_vectors_ready,
      BatchIn_vectors_dvalid        => Abs_kernel_Nucleus_inst_BatchIn_vectors_dvalid,
      BatchIn_vectors_last          => Abs_kernel_Nucleus_inst_BatchIn_vectors_last,
      BatchIn_vectors               => Abs_kernel_Nucleus_inst_BatchIn_vectors,
      BatchIn_vectors_unl_valid     => Abs_kernel_Nucleus_inst_BatchIn_vectors_unl_valid,
      BatchIn_vectors_unl_ready     => Abs_kernel_Nucleus_inst_BatchIn_vectors_unl_ready,
      BatchIn_vectors_unl_tag       => Abs_kernel_Nucleus_inst_BatchIn_vectors_unl_tag,
      BatchIn_vectors_cmd_valid     => Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_valid,
      BatchIn_vectors_cmd_ready     => Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_ready,
      BatchIn_vectors_cmd_firstIdx  => Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_firstIdx,
      BatchIn_vectors_cmd_lastIdx   => Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_lastIdx,
      BatchIn_vectors_cmd_ctrl      => Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_ctrl,
      BatchIn_vectors_cmd_tag       => Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_tag,
      BatchOut_vectors_valid        => Abs_kernel_Nucleus_inst_BatchOut_vectors_valid,
      BatchOut_vectors_ready        => Abs_kernel_Nucleus_inst_BatchOut_vectors_ready,
      BatchOut_vectors_dvalid       => Abs_kernel_Nucleus_inst_BatchOut_vectors_dvalid,
      BatchOut_vectors_last         => Abs_kernel_Nucleus_inst_BatchOut_vectors_last,
      BatchOut_vectors              => Abs_kernel_Nucleus_inst_BatchOut_vectors,
      BatchOut_vectors_unl_valid    => Abs_kernel_Nucleus_inst_BatchOut_vectors_unl_valid,
      BatchOut_vectors_unl_ready    => Abs_kernel_Nucleus_inst_BatchOut_vectors_unl_ready,
      BatchOut_vectors_unl_tag      => Abs_kernel_Nucleus_inst_BatchOut_vectors_unl_tag,
      BatchOut_vectors_cmd_valid    => Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_valid,
      BatchOut_vectors_cmd_ready    => Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_ready,
      BatchOut_vectors_cmd_firstIdx => Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_firstIdx,
      BatchOut_vectors_cmd_lastIdx  => Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_lastIdx,
      BatchOut_vectors_cmd_ctrl     => Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_ctrl,
      BatchOut_vectors_cmd_tag      => Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_tag
    );

  Abs_kernel_BatchIn_inst : Abs_kernel_BatchIn
    generic map (
      INDEX_WIDTH                        => INDEX_WIDTH,
      TAG_WIDTH                          => TAG_WIDTH,
      BATCHIN_VECTORS_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      BATCHIN_VECTORS_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      BATCHIN_VECTORS_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      BATCHIN_VECTORS_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      BATCHIN_VECTORS_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                        => Abs_kernel_BatchIn_inst_bcd_clk,
      bcd_reset                      => Abs_kernel_BatchIn_inst_bcd_reset,
      kcd_clk                        => Abs_kernel_BatchIn_inst_kcd_clk,
      kcd_reset                      => Abs_kernel_BatchIn_inst_kcd_reset,
      BatchIn_vectors_valid          => Abs_kernel_BatchIn_inst_BatchIn_vectors_valid,
      BatchIn_vectors_ready          => Abs_kernel_BatchIn_inst_BatchIn_vectors_ready,
      BatchIn_vectors_dvalid         => Abs_kernel_BatchIn_inst_BatchIn_vectors_dvalid,
      BatchIn_vectors_last           => Abs_kernel_BatchIn_inst_BatchIn_vectors_last,
      BatchIn_vectors                => Abs_kernel_BatchIn_inst_BatchIn_vectors,
      BatchIn_vectors_bus_rreq_valid => Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rreq_valid,
      BatchIn_vectors_bus_rreq_ready => Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rreq_ready,
      BatchIn_vectors_bus_rreq_addr  => Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rreq_addr,
      BatchIn_vectors_bus_rreq_len   => Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rreq_len,
      BatchIn_vectors_bus_rdat_valid => Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rdat_valid,
      BatchIn_vectors_bus_rdat_ready => Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rdat_ready,
      BatchIn_vectors_bus_rdat_data  => Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rdat_data,
      BatchIn_vectors_bus_rdat_last  => Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rdat_last,
      BatchIn_vectors_cmd_valid      => Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_valid,
      BatchIn_vectors_cmd_ready      => Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_ready,
      BatchIn_vectors_cmd_firstIdx   => Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_firstIdx,
      BatchIn_vectors_cmd_lastIdx    => Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_lastIdx,
      BatchIn_vectors_cmd_ctrl       => Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_ctrl,
      BatchIn_vectors_cmd_tag        => Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_tag,
      BatchIn_vectors_unl_valid      => Abs_kernel_BatchIn_inst_BatchIn_vectors_unl_valid,
      BatchIn_vectors_unl_ready      => Abs_kernel_BatchIn_inst_BatchIn_vectors_unl_ready,
      BatchIn_vectors_unl_tag        => Abs_kernel_BatchIn_inst_BatchIn_vectors_unl_tag
    );

  Abs_kernel_BatchOut_inst : Abs_kernel_BatchOut
    generic map (
      INDEX_WIDTH                         => INDEX_WIDTH,
      TAG_WIDTH                           => TAG_WIDTH,
      BATCHOUT_VECTORS_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      BATCHOUT_VECTORS_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      BATCHOUT_VECTORS_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      BATCHOUT_VECTORS_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      BATCHOUT_VECTORS_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                          => Abs_kernel_BatchOut_inst_bcd_clk,
      bcd_reset                        => Abs_kernel_BatchOut_inst_bcd_reset,
      kcd_clk                          => Abs_kernel_BatchOut_inst_kcd_clk,
      kcd_reset                        => Abs_kernel_BatchOut_inst_kcd_reset,
      BatchOut_vectors_valid           => Abs_kernel_BatchOut_inst_BatchOut_vectors_valid,
      BatchOut_vectors_ready           => Abs_kernel_BatchOut_inst_BatchOut_vectors_ready,
      BatchOut_vectors_dvalid          => Abs_kernel_BatchOut_inst_BatchOut_vectors_dvalid,
      BatchOut_vectors_last            => Abs_kernel_BatchOut_inst_BatchOut_vectors_last,
      BatchOut_vectors                 => Abs_kernel_BatchOut_inst_BatchOut_vectors,
      BatchOut_vectors_bus_wreq_valid  => Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wreq_valid,
      BatchOut_vectors_bus_wreq_ready  => Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wreq_ready,
      BatchOut_vectors_bus_wreq_addr   => Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wreq_addr,
      BatchOut_vectors_bus_wreq_len    => Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wreq_len,
      BatchOut_vectors_bus_wdat_valid  => Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_valid,
      BatchOut_vectors_bus_wdat_ready  => Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_ready,
      BatchOut_vectors_bus_wdat_data   => Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_data,
      BatchOut_vectors_bus_wdat_strobe => Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_strobe,
      BatchOut_vectors_bus_wdat_last   => Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_last,
      BatchOut_vectors_cmd_valid       => Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_valid,
      BatchOut_vectors_cmd_ready       => Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_ready,
      BatchOut_vectors_cmd_firstIdx    => Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_firstIdx,
      BatchOut_vectors_cmd_lastIdx     => Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_lastIdx,
      BatchOut_vectors_cmd_ctrl        => Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_ctrl,
      BatchOut_vectors_cmd_tag         => Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_tag,
      BatchOut_vectors_unl_valid       => Abs_kernel_BatchOut_inst_BatchOut_vectors_unl_valid,
      BatchOut_vectors_unl_ready       => Abs_kernel_BatchOut_inst_BatchOut_vectors_unl_ready,
      BatchOut_vectors_unl_tag         => Abs_kernel_BatchOut_inst_BatchOut_vectors_unl_tag
    );

  RDAW64DW512LW8BS1BM16_inst : BusReadArbiterVec
    generic map (
      BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH  => BUS_DATA_WIDTH,
      BUS_LEN_WIDTH   => BUS_LEN_WIDTH,
      NUM_SLAVE_PORTS => 1,
      ARB_METHOD      => "RR-STICKY",
      MAX_OUTSTANDING => 4,
      RAM_CONFIG      => "",
      SLV_REQ_SLICES  => true,
      MST_REQ_SLICE   => true,
      MST_DAT_SLICE   => true,
      SLV_DAT_SLICES  => true
    )
    port map (
      bcd_clk        => RDAW64DW512LW8BS1BM16_inst_bcd_clk,
      bcd_reset      => RDAW64DW512LW8BS1BM16_inst_bcd_reset,
      mst_rreq_valid => RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid,
      mst_rreq_ready => RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready,
      mst_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr,
      mst_rreq_len   => RDAW64DW512LW8BS1BM16_inst_mst_rreq_len,
      mst_rdat_valid => RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid,
      mst_rdat_ready => RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready,
      mst_rdat_data  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_data,
      mst_rdat_last  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_last,
      bsv_rreq_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid,
      bsv_rreq_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready,
      bsv_rreq_len   => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len,
      bsv_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr,
      bsv_rdat_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid,
      bsv_rdat_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready,
      bsv_rdat_last  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last,
      bsv_rdat_data  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data
    );

  WRAW64DW512LW8BS1BM16_inst : BusWriteArbiterVec
    generic map (
      BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH  => BUS_DATA_WIDTH,
      BUS_LEN_WIDTH   => BUS_LEN_WIDTH,
      NUM_SLAVE_PORTS => 1,
      ARB_METHOD      => "RR-STICKY",
      MAX_OUTSTANDING => 4,
      RAM_CONFIG      => "",
      SLV_REQ_SLICES  => true,
      MST_REQ_SLICE   => true,
      MST_DAT_SLICE   => true,
      SLV_DAT_SLICES  => true
    )
    port map (
      bcd_clk         => WRAW64DW512LW8BS1BM16_inst_bcd_clk,
      bcd_reset       => WRAW64DW512LW8BS1BM16_inst_bcd_reset,
      mst_wreq_valid  => WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid,
      mst_wreq_ready  => WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready,
      mst_wreq_addr   => WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr,
      mst_wreq_len    => WRAW64DW512LW8BS1BM16_inst_mst_wreq_len,
      mst_wdat_valid  => WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid,
      mst_wdat_ready  => WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready,
      mst_wdat_data   => WRAW64DW512LW8BS1BM16_inst_mst_wdat_data,
      mst_wdat_strobe => WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe,
      mst_wdat_last   => WRAW64DW512LW8BS1BM16_inst_mst_wdat_last,
      bsv_wreq_valid  => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid,
      bsv_wreq_ready  => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready,
      bsv_wreq_len    => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len,
      bsv_wreq_addr   => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr,
      bsv_wdat_valid  => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid,
      bsv_wdat_strobe => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe,
      bsv_wdat_ready  => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready,
      bsv_wdat_last   => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last,
      bsv_wdat_data   => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data
    );

  rd_mst_rreq_valid                         <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready <= rd_mst_rreq_ready;
  rd_mst_rreq_addr                          <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr;
  rd_mst_rreq_len                           <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid <= rd_mst_rdat_valid;
  rd_mst_rdat_ready                         <= RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_data  <= rd_mst_rdat_data;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_last  <= rd_mst_rdat_last;

  wr_mst_wreq_valid                         <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready <= wr_mst_wreq_ready;
  wr_mst_wreq_addr                          <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr;
  wr_mst_wreq_len                           <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_len;
  wr_mst_wdat_valid                         <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready <= wr_mst_wdat_ready;
  wr_mst_wdat_data                          <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_data;
  wr_mst_wdat_strobe                        <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe;
  wr_mst_wdat_last                          <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_last;

  Abs_kernel_Nucleus_inst_kcd_clk                        <= kcd_clk;
  Abs_kernel_Nucleus_inst_kcd_reset                      <= kcd_reset;

  Abs_kernel_Nucleus_inst_mmio_awvalid                   <= mmio_awvalid;
  mmio_awready                                           <= Abs_kernel_Nucleus_inst_mmio_awready;
  Abs_kernel_Nucleus_inst_mmio_awaddr                    <= mmio_awaddr;
  Abs_kernel_Nucleus_inst_mmio_wvalid                    <= mmio_wvalid;
  mmio_wready                                            <= Abs_kernel_Nucleus_inst_mmio_wready;
  Abs_kernel_Nucleus_inst_mmio_wdata                     <= mmio_wdata;
  Abs_kernel_Nucleus_inst_mmio_wstrb                     <= mmio_wstrb;
  mmio_bvalid                                            <= Abs_kernel_Nucleus_inst_mmio_bvalid;
  Abs_kernel_Nucleus_inst_mmio_bready                    <= mmio_bready;
  mmio_bresp                                             <= Abs_kernel_Nucleus_inst_mmio_bresp;
  Abs_kernel_Nucleus_inst_mmio_arvalid                   <= mmio_arvalid;
  mmio_arready                                           <= Abs_kernel_Nucleus_inst_mmio_arready;
  Abs_kernel_Nucleus_inst_mmio_araddr                    <= mmio_araddr;
  mmio_rvalid                                            <= Abs_kernel_Nucleus_inst_mmio_rvalid;
  Abs_kernel_Nucleus_inst_mmio_rready                    <= mmio_rready;
  mmio_rdata                                             <= Abs_kernel_Nucleus_inst_mmio_rdata;
  mmio_rresp                                             <= Abs_kernel_Nucleus_inst_mmio_rresp;

  Abs_kernel_Nucleus_inst_BatchIn_vectors_valid          <= Abs_kernel_BatchIn_inst_BatchIn_vectors_valid;
  Abs_kernel_BatchIn_inst_BatchIn_vectors_ready          <= Abs_kernel_Nucleus_inst_BatchIn_vectors_ready;
  Abs_kernel_Nucleus_inst_BatchIn_vectors_dvalid         <= Abs_kernel_BatchIn_inst_BatchIn_vectors_dvalid;
  Abs_kernel_Nucleus_inst_BatchIn_vectors_last           <= Abs_kernel_BatchIn_inst_BatchIn_vectors_last;
  Abs_kernel_Nucleus_inst_BatchIn_vectors                <= Abs_kernel_BatchIn_inst_BatchIn_vectors;

  Abs_kernel_Nucleus_inst_BatchIn_vectors_unl_valid      <= Abs_kernel_BatchIn_inst_BatchIn_vectors_unl_valid;
  Abs_kernel_BatchIn_inst_BatchIn_vectors_unl_ready      <= Abs_kernel_Nucleus_inst_BatchIn_vectors_unl_ready;
  Abs_kernel_Nucleus_inst_BatchIn_vectors_unl_tag        <= Abs_kernel_BatchIn_inst_BatchIn_vectors_unl_tag;

  Abs_kernel_Nucleus_inst_BatchOut_vectors_unl_valid     <= Abs_kernel_BatchOut_inst_BatchOut_vectors_unl_valid;
  Abs_kernel_BatchOut_inst_BatchOut_vectors_unl_ready    <= Abs_kernel_Nucleus_inst_BatchOut_vectors_unl_ready;
  Abs_kernel_Nucleus_inst_BatchOut_vectors_unl_tag       <= Abs_kernel_BatchOut_inst_BatchOut_vectors_unl_tag;

  Abs_kernel_BatchIn_inst_bcd_clk                        <= bcd_clk;
  Abs_kernel_BatchIn_inst_bcd_reset                      <= bcd_reset;

  Abs_kernel_BatchIn_inst_kcd_clk                        <= kcd_clk;
  Abs_kernel_BatchIn_inst_kcd_reset                      <= kcd_reset;

  Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_valid      <= Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_valid;
  Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_ready      <= Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_ready;
  Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_firstIdx   <= Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_firstIdx;
  Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_lastIdx    <= Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_lastIdx;
  Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_ctrl       <= Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_ctrl;
  Abs_kernel_BatchIn_inst_BatchIn_vectors_cmd_tag        <= Abs_kernel_Nucleus_inst_BatchIn_vectors_cmd_tag;

  Abs_kernel_BatchOut_inst_bcd_clk                       <= bcd_clk;
  Abs_kernel_BatchOut_inst_bcd_reset                     <= bcd_reset;

  Abs_kernel_BatchOut_inst_kcd_clk                       <= kcd_clk;
  Abs_kernel_BatchOut_inst_kcd_reset                     <= kcd_reset;

  Abs_kernel_BatchOut_inst_BatchOut_vectors_valid        <= Abs_kernel_Nucleus_inst_BatchOut_vectors_valid;
  Abs_kernel_Nucleus_inst_BatchOut_vectors_ready         <= Abs_kernel_BatchOut_inst_BatchOut_vectors_ready;
  Abs_kernel_BatchOut_inst_BatchOut_vectors_dvalid       <= Abs_kernel_Nucleus_inst_BatchOut_vectors_dvalid;
  Abs_kernel_BatchOut_inst_BatchOut_vectors_last         <= Abs_kernel_Nucleus_inst_BatchOut_vectors_last;
  Abs_kernel_BatchOut_inst_BatchOut_vectors              <= Abs_kernel_Nucleus_inst_BatchOut_vectors;

  Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_valid    <= Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_valid;
  Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_ready     <= Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_ready;
  Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_firstIdx <= Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_firstIdx;
  Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_lastIdx  <= Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_lastIdx;
  Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_ctrl     <= Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_ctrl;
  Abs_kernel_BatchOut_inst_BatchOut_vectors_cmd_tag      <= Abs_kernel_Nucleus_inst_BatchOut_vectors_cmd_tag;

  RDAW64DW512LW8BS1BM16_inst_bcd_clk                     <= bcd_clk;
  RDAW64DW512LW8BS1BM16_inst_bcd_reset                   <= bcd_reset;

  WRAW64DW512LW8BS1BM16_inst_bcd_clk                     <= bcd_clk;
  WRAW64DW512LW8BS1BM16_inst_bcd_reset                   <= bcd_reset;

  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(0)                            <= Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH-1 downto 0)       <= Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH-1 downto 0)     <= Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(0)                            <= Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rdat_ready;
  Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rreq_ready                  <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(0);
  Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rdat_valid                  <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(0);
  Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rdat_last                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(0);
  Abs_kernel_BatchIn_inst_BatchIn_vectors_bus_rdat_data                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH-1 downto 0);

  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(0)                            <= Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH-1 downto 0)       <= Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH-1 downto 0)     <= Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(0)                            <= Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8-1 downto 0) <= Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(0)                             <= Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH-1 downto 0)     <= Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_data;
  Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wreq_ready                <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(0);
  Abs_kernel_BatchOut_inst_BatchOut_vectors_bus_wdat_ready                <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(0);

end architecture;
