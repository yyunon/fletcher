-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;

entity Abs_kernel_BatchIn is
  generic (
    INDEX_WIDTH                        : integer := 32;
    TAG_WIDTH                          : integer := 1;
    BATCHIN_VECTORS_BUS_ADDR_WIDTH     : integer := 64;
    BATCHIN_VECTORS_BUS_DATA_WIDTH     : integer := 512;
    BATCHIN_VECTORS_BUS_LEN_WIDTH      : integer := 8;
    BATCHIN_VECTORS_BUS_BURST_STEP_LEN : integer := 1;
    BATCHIN_VECTORS_BUS_BURST_MAX_LEN  : integer := 16
  );
  port (
    bcd_clk                        : in  std_logic;
    bcd_reset                      : in  std_logic;
    kcd_clk                        : in  std_logic;
    kcd_reset                      : in  std_logic;
    BatchIn_vectors_valid          : out std_logic;
    BatchIn_vectors_ready          : in  std_logic;
    BatchIn_vectors_dvalid         : out std_logic;
    BatchIn_vectors_last           : out std_logic;
    BatchIn_vectors                : out std_logic_vector(63 downto 0);
    BatchIn_vectors_bus_rreq_valid : out std_logic;
    BatchIn_vectors_bus_rreq_ready : in  std_logic;
    BatchIn_vectors_bus_rreq_addr  : out std_logic_vector(BATCHIN_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
    BatchIn_vectors_bus_rreq_len   : out std_logic_vector(BATCHIN_VECTORS_BUS_LEN_WIDTH-1 downto 0);
    BatchIn_vectors_bus_rdat_valid : in  std_logic;
    BatchIn_vectors_bus_rdat_ready : out std_logic;
    BatchIn_vectors_bus_rdat_data  : in  std_logic_vector(BATCHIN_VECTORS_BUS_DATA_WIDTH-1 downto 0);
    BatchIn_vectors_bus_rdat_last  : in  std_logic;
    BatchIn_vectors_cmd_valid      : in  std_logic;
    BatchIn_vectors_cmd_ready      : out std_logic;
    BatchIn_vectors_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    BatchIn_vectors_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    BatchIn_vectors_cmd_ctrl       : in  std_logic_vector(BATCHIN_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
    BatchIn_vectors_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    BatchIn_vectors_unl_valid      : out std_logic;
    BatchIn_vectors_unl_ready      : in  std_logic;
    BatchIn_vectors_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
  );
end entity;

architecture Implementation of Abs_kernel_BatchIn is
  signal vectors_inst_bcd_clk        : std_logic;
  signal vectors_inst_bcd_reset      : std_logic;

  signal vectors_inst_kcd_clk        : std_logic;
  signal vectors_inst_kcd_reset      : std_logic;

  signal vectors_inst_cmd_valid      : std_logic;
  signal vectors_inst_cmd_ready      : std_logic;
  signal vectors_inst_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal vectors_inst_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal vectors_inst_cmd_ctrl       : std_logic_vector(BATCHIN_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
  signal vectors_inst_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal vectors_inst_unl_valid      : std_logic;
  signal vectors_inst_unl_ready      : std_logic;
  signal vectors_inst_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal vectors_inst_bus_rreq_valid : std_logic;
  signal vectors_inst_bus_rreq_ready : std_logic;
  signal vectors_inst_bus_rreq_addr  : std_logic_vector(BATCHIN_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
  signal vectors_inst_bus_rreq_len   : std_logic_vector(BATCHIN_VECTORS_BUS_LEN_WIDTH-1 downto 0);
  signal vectors_inst_bus_rdat_valid : std_logic;
  signal vectors_inst_bus_rdat_ready : std_logic;
  signal vectors_inst_bus_rdat_data  : std_logic_vector(BATCHIN_VECTORS_BUS_DATA_WIDTH-1 downto 0);
  signal vectors_inst_bus_rdat_last  : std_logic;

  signal vectors_inst_out_valid      : std_logic_vector(0 downto 0);
  signal vectors_inst_out_ready      : std_logic_vector(0 downto 0);
  signal vectors_inst_out_data       : std_logic_vector(63 downto 0);
  signal vectors_inst_out_dvalid     : std_logic_vector(0 downto 0);
  signal vectors_inst_out_last       : std_logic_vector(0 downto 0);

begin
  vectors_inst : ArrayReader
    generic map (
      BUS_ADDR_WIDTH     => BATCHIN_VECTORS_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => BATCHIN_VECTORS_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => BATCHIN_VECTORS_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => BATCHIN_VECTORS_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => BATCHIN_VECTORS_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk        => vectors_inst_bcd_clk,
      bcd_reset      => vectors_inst_bcd_reset,
      kcd_clk        => vectors_inst_kcd_clk,
      kcd_reset      => vectors_inst_kcd_reset,
      cmd_valid      => vectors_inst_cmd_valid,
      cmd_ready      => vectors_inst_cmd_ready,
      cmd_firstIdx   => vectors_inst_cmd_firstIdx,
      cmd_lastIdx    => vectors_inst_cmd_lastIdx,
      cmd_ctrl       => vectors_inst_cmd_ctrl,
      cmd_tag        => vectors_inst_cmd_tag,
      unl_valid      => vectors_inst_unl_valid,
      unl_ready      => vectors_inst_unl_ready,
      unl_tag        => vectors_inst_unl_tag,
      bus_rreq_valid => vectors_inst_bus_rreq_valid,
      bus_rreq_ready => vectors_inst_bus_rreq_ready,
      bus_rreq_addr  => vectors_inst_bus_rreq_addr,
      bus_rreq_len   => vectors_inst_bus_rreq_len,
      bus_rdat_valid => vectors_inst_bus_rdat_valid,
      bus_rdat_ready => vectors_inst_bus_rdat_ready,
      bus_rdat_data  => vectors_inst_bus_rdat_data,
      bus_rdat_last  => vectors_inst_bus_rdat_last,
      out_valid      => vectors_inst_out_valid,
      out_ready      => vectors_inst_out_ready,
      out_data       => vectors_inst_out_data,
      out_dvalid     => vectors_inst_out_dvalid,
      out_last       => vectors_inst_out_last
    );

  BatchIn_vectors_valid          <= vectors_inst_out_valid(0);
  vectors_inst_out_ready(0)      <= BatchIn_vectors_ready;
  BatchIn_vectors_dvalid         <= vectors_inst_out_dvalid(0);
  BatchIn_vectors_last           <= vectors_inst_out_last(0);
  BatchIn_vectors                <= vectors_inst_out_data;

  BatchIn_vectors_bus_rreq_valid <= vectors_inst_bus_rreq_valid;
  vectors_inst_bus_rreq_ready    <= BatchIn_vectors_bus_rreq_ready;
  BatchIn_vectors_bus_rreq_addr  <= vectors_inst_bus_rreq_addr;
  BatchIn_vectors_bus_rreq_len   <= vectors_inst_bus_rreq_len;
  vectors_inst_bus_rdat_valid    <= BatchIn_vectors_bus_rdat_valid;
  BatchIn_vectors_bus_rdat_ready <= vectors_inst_bus_rdat_ready;
  vectors_inst_bus_rdat_data     <= BatchIn_vectors_bus_rdat_data;
  vectors_inst_bus_rdat_last     <= BatchIn_vectors_bus_rdat_last;

  BatchIn_vectors_unl_valid      <= vectors_inst_unl_valid;
  vectors_inst_unl_ready         <= BatchIn_vectors_unl_ready;
  BatchIn_vectors_unl_tag        <= vectors_inst_unl_tag;

  vectors_inst_bcd_clk      <= bcd_clk;
  vectors_inst_bcd_reset    <= bcd_reset;

  vectors_inst_kcd_clk      <= kcd_clk;
  vectors_inst_kcd_reset    <= kcd_reset;

  vectors_inst_cmd_valid    <= BatchIn_vectors_cmd_valid;
  BatchIn_vectors_cmd_ready <= vectors_inst_cmd_ready;
  vectors_inst_cmd_firstIdx <= BatchIn_vectors_cmd_firstIdx;
  vectors_inst_cmd_lastIdx  <= BatchIn_vectors_cmd_lastIdx;
  vectors_inst_cmd_ctrl     <= BatchIn_vectors_cmd_ctrl;
  vectors_inst_cmd_tag      <= BatchIn_vectors_cmd_tag;

end architecture;
