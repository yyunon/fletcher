-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Interconnect_pkg.all;

entity Sum_Mantle is
  generic (
    INDEX_WIDTH        : integer := 32;
    TAG_WIDTH          : integer := 1;
    BUS_ADDR_WIDTH     : integer := 64;
    BUS_DATA_WIDTH     : integer := 512;
    BUS_LEN_WIDTH      : integer := 8;
    BUS_BURST_STEP_LEN : integer := 1;
    BUS_BURST_MAX_LEN  : integer := 16
  );
  port (
    bcd_clk           : in  std_logic;
    bcd_reset         : in  std_logic;
    kcd_clk           : in  std_logic;
    kcd_reset         : in  std_logic;
    mmio_awvalid      : in  std_logic;
    mmio_awready      : out std_logic;
    mmio_awaddr       : in  std_logic_vector(31 downto 0);
    mmio_wvalid       : in  std_logic;
    mmio_wready       : out std_logic;
    mmio_wdata        : in  std_logic_vector(31 downto 0);
    mmio_wstrb        : in  std_logic_vector(3 downto 0);
    mmio_bvalid       : out std_logic;
    mmio_bready       : in  std_logic;
    mmio_bresp        : out std_logic_vector(1 downto 0);
    mmio_arvalid      : in  std_logic;
    mmio_arready      : out std_logic;
    mmio_araddr       : in  std_logic_vector(31 downto 0);
    mmio_rvalid       : out std_logic;
    mmio_rready       : in  std_logic;
    mmio_rdata        : out std_logic_vector(31 downto 0);
    mmio_rresp        : out std_logic_vector(1 downto 0);
    rd_mst_rreq_valid : out std_logic;
    rd_mst_rreq_ready : in  std_logic;
    rd_mst_rreq_addr  : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    rd_mst_rreq_len   : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    rd_mst_rdat_valid : in  std_logic;
    rd_mst_rdat_ready : out std_logic;
    rd_mst_rdat_data  : in  std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    rd_mst_rdat_last  : in  std_logic
  );
end entity;

architecture Implementation of Sum_Mantle is
  component Sum_Nucleus is
    generic (
      INDEX_WIDTH                        : integer := 32;
      TAG_WIDTH                          : integer := 1;
      EXAMPLEBATCH_NUMBER_BUS_ADDR_WIDTH : integer := 64
    );
    port (
      kcd_clk                          : in  std_logic;
      kcd_reset                        : in  std_logic;
      mmio_awvalid                     : in  std_logic;
      mmio_awready                     : out std_logic;
      mmio_awaddr                      : in  std_logic_vector(31 downto 0);
      mmio_wvalid                      : in  std_logic;
      mmio_wready                      : out std_logic;
      mmio_wdata                       : in  std_logic_vector(31 downto 0);
      mmio_wstrb                       : in  std_logic_vector(3 downto 0);
      mmio_bvalid                      : out std_logic;
      mmio_bready                      : in  std_logic;
      mmio_bresp                       : out std_logic_vector(1 downto 0);
      mmio_arvalid                     : in  std_logic;
      mmio_arready                     : out std_logic;
      mmio_araddr                      : in  std_logic_vector(31 downto 0);
      mmio_rvalid                      : out std_logic;
      mmio_rready                      : in  std_logic;
      mmio_rdata                       : out std_logic_vector(31 downto 0);
      mmio_rresp                       : out std_logic_vector(1 downto 0);
      ExampleBatch_number_valid        : in  std_logic;
      ExampleBatch_number_ready        : out std_logic;
      ExampleBatch_number_dvalid       : in  std_logic;
      ExampleBatch_number_last         : in  std_logic;
      ExampleBatch_number              : in  std_logic_vector(63 downto 0);
      ExampleBatch_number_unl_valid    : in  std_logic;
      ExampleBatch_number_unl_ready    : out std_logic;
      ExampleBatch_number_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ExampleBatch_number_cmd_valid    : out std_logic;
      ExampleBatch_number_cmd_ready    : in  std_logic;
      ExampleBatch_number_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ExampleBatch_number_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ExampleBatch_number_cmd_ctrl     : out std_logic_vector(EXAMPLEBATCH_NUMBER_BUS_ADDR_WIDTH-1 downto 0);
      ExampleBatch_number_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Sum_ExampleBatch is
    generic (
      INDEX_WIDTH                            : integer := 32;
      TAG_WIDTH                              : integer := 1;
      EXAMPLEBATCH_NUMBER_BUS_ADDR_WIDTH     : integer := 64;
      EXAMPLEBATCH_NUMBER_BUS_DATA_WIDTH     : integer := 512;
      EXAMPLEBATCH_NUMBER_BUS_LEN_WIDTH      : integer := 8;
      EXAMPLEBATCH_NUMBER_BUS_BURST_STEP_LEN : integer := 1;
      EXAMPLEBATCH_NUMBER_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                            : in  std_logic;
      bcd_reset                          : in  std_logic;
      kcd_clk                            : in  std_logic;
      kcd_reset                          : in  std_logic;
      ExampleBatch_number_valid          : out std_logic;
      ExampleBatch_number_ready          : in  std_logic;
      ExampleBatch_number_dvalid         : out std_logic;
      ExampleBatch_number_last           : out std_logic;
      ExampleBatch_number                : out std_logic_vector(63 downto 0);
      ExampleBatch_number_bus_rreq_valid : out std_logic;
      ExampleBatch_number_bus_rreq_ready : in  std_logic;
      ExampleBatch_number_bus_rreq_addr  : out std_logic_vector(EXAMPLEBATCH_NUMBER_BUS_ADDR_WIDTH-1 downto 0);
      ExampleBatch_number_bus_rreq_len   : out std_logic_vector(EXAMPLEBATCH_NUMBER_BUS_LEN_WIDTH-1 downto 0);
      ExampleBatch_number_bus_rdat_valid : in  std_logic;
      ExampleBatch_number_bus_rdat_ready : out std_logic;
      ExampleBatch_number_bus_rdat_data  : in  std_logic_vector(EXAMPLEBATCH_NUMBER_BUS_DATA_WIDTH-1 downto 0);
      ExampleBatch_number_bus_rdat_last  : in  std_logic;
      ExampleBatch_number_cmd_valid      : in  std_logic;
      ExampleBatch_number_cmd_ready      : out std_logic;
      ExampleBatch_number_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ExampleBatch_number_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ExampleBatch_number_cmd_ctrl       : in  std_logic_vector(EXAMPLEBATCH_NUMBER_BUS_ADDR_WIDTH-1 downto 0);
      ExampleBatch_number_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ExampleBatch_number_unl_valid      : out std_logic;
      ExampleBatch_number_unl_ready      : in  std_logic;
      ExampleBatch_number_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  signal Sum_Nucleus_inst_kcd_clk                                 : std_logic;
  signal Sum_Nucleus_inst_kcd_reset                               : std_logic;

  signal Sum_Nucleus_inst_mmio_awvalid                            : std_logic;
  signal Sum_Nucleus_inst_mmio_awready                            : std_logic;
  signal Sum_Nucleus_inst_mmio_awaddr                             : std_logic_vector(31 downto 0);
  signal Sum_Nucleus_inst_mmio_wvalid                             : std_logic;
  signal Sum_Nucleus_inst_mmio_wready                             : std_logic;
  signal Sum_Nucleus_inst_mmio_wdata                              : std_logic_vector(31 downto 0);
  signal Sum_Nucleus_inst_mmio_wstrb                              : std_logic_vector(3 downto 0);
  signal Sum_Nucleus_inst_mmio_bvalid                             : std_logic;
  signal Sum_Nucleus_inst_mmio_bready                             : std_logic;
  signal Sum_Nucleus_inst_mmio_bresp                              : std_logic_vector(1 downto 0);
  signal Sum_Nucleus_inst_mmio_arvalid                            : std_logic;
  signal Sum_Nucleus_inst_mmio_arready                            : std_logic;
  signal Sum_Nucleus_inst_mmio_araddr                             : std_logic_vector(31 downto 0);
  signal Sum_Nucleus_inst_mmio_rvalid                             : std_logic;
  signal Sum_Nucleus_inst_mmio_rready                             : std_logic;
  signal Sum_Nucleus_inst_mmio_rdata                              : std_logic_vector(31 downto 0);
  signal Sum_Nucleus_inst_mmio_rresp                              : std_logic_vector(1 downto 0);

  signal Sum_Nucleus_inst_ExampleBatch_number_valid               : std_logic;
  signal Sum_Nucleus_inst_ExampleBatch_number_ready               : std_logic;
  signal Sum_Nucleus_inst_ExampleBatch_number_dvalid              : std_logic;
  signal Sum_Nucleus_inst_ExampleBatch_number_last                : std_logic;
  signal Sum_Nucleus_inst_ExampleBatch_number                     : std_logic_vector(63 downto 0);

  signal Sum_Nucleus_inst_ExampleBatch_number_unl_valid           : std_logic;
  signal Sum_Nucleus_inst_ExampleBatch_number_unl_ready           : std_logic;
  signal Sum_Nucleus_inst_ExampleBatch_number_unl_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Sum_Nucleus_inst_ExampleBatch_number_cmd_valid           : std_logic;
  signal Sum_Nucleus_inst_ExampleBatch_number_cmd_ready           : std_logic;
  signal Sum_Nucleus_inst_ExampleBatch_number_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Sum_Nucleus_inst_ExampleBatch_number_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Sum_Nucleus_inst_ExampleBatch_number_cmd_ctrl            : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Sum_Nucleus_inst_ExampleBatch_number_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Sum_ExampleBatch_inst_bcd_clk                            : std_logic;
  signal Sum_ExampleBatch_inst_bcd_reset                          : std_logic;

  signal Sum_ExampleBatch_inst_kcd_clk                            : std_logic;
  signal Sum_ExampleBatch_inst_kcd_reset                          : std_logic;

  signal Sum_ExampleBatch_inst_ExampleBatch_number_valid          : std_logic;
  signal Sum_ExampleBatch_inst_ExampleBatch_number_ready          : std_logic;
  signal Sum_ExampleBatch_inst_ExampleBatch_number_dvalid         : std_logic;
  signal Sum_ExampleBatch_inst_ExampleBatch_number_last           : std_logic;
  signal Sum_ExampleBatch_inst_ExampleBatch_number                : std_logic_vector(63 downto 0);

  signal Sum_ExampleBatch_inst_ExampleBatch_number_bus_rreq_valid : std_logic;
  signal Sum_ExampleBatch_inst_ExampleBatch_number_bus_rreq_ready : std_logic;
  signal Sum_ExampleBatch_inst_ExampleBatch_number_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Sum_ExampleBatch_inst_ExampleBatch_number_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Sum_ExampleBatch_inst_ExampleBatch_number_bus_rdat_valid : std_logic;
  signal Sum_ExampleBatch_inst_ExampleBatch_number_bus_rdat_ready : std_logic;
  signal Sum_ExampleBatch_inst_ExampleBatch_number_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Sum_ExampleBatch_inst_ExampleBatch_number_bus_rdat_last  : std_logic;

  signal Sum_ExampleBatch_inst_ExampleBatch_number_cmd_valid      : std_logic;
  signal Sum_ExampleBatch_inst_ExampleBatch_number_cmd_ready      : std_logic;
  signal Sum_ExampleBatch_inst_ExampleBatch_number_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Sum_ExampleBatch_inst_ExampleBatch_number_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Sum_ExampleBatch_inst_ExampleBatch_number_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Sum_ExampleBatch_inst_ExampleBatch_number_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Sum_ExampleBatch_inst_ExampleBatch_number_unl_valid      : std_logic;
  signal Sum_ExampleBatch_inst_ExampleBatch_number_unl_ready      : std_logic;
  signal Sum_ExampleBatch_inst_ExampleBatch_number_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal RDAW64DW512LW8BS1BM16_inst_bcd_clk                       : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_bcd_reset                     : std_logic;

  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid                : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready                : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr                 : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_len                  : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid                : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready                : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_data                 : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_last                 : std_logic;

  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid : std_logic_vector(0 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready : std_logic_vector(0 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid : std_logic_vector(0 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready : std_logic_vector(0 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last  : std_logic_vector(0 downto 0);

begin
  Sum_Nucleus_inst : Sum_Nucleus
    generic map (
      INDEX_WIDTH                        => INDEX_WIDTH,
      TAG_WIDTH                          => TAG_WIDTH,
      EXAMPLEBATCH_NUMBER_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH
    )
    port map (
      kcd_clk                          => Sum_Nucleus_inst_kcd_clk,
      kcd_reset                        => Sum_Nucleus_inst_kcd_reset,
      mmio_awvalid                     => Sum_Nucleus_inst_mmio_awvalid,
      mmio_awready                     => Sum_Nucleus_inst_mmio_awready,
      mmio_awaddr                      => Sum_Nucleus_inst_mmio_awaddr,
      mmio_wvalid                      => Sum_Nucleus_inst_mmio_wvalid,
      mmio_wready                      => Sum_Nucleus_inst_mmio_wready,
      mmio_wdata                       => Sum_Nucleus_inst_mmio_wdata,
      mmio_wstrb                       => Sum_Nucleus_inst_mmio_wstrb,
      mmio_bvalid                      => Sum_Nucleus_inst_mmio_bvalid,
      mmio_bready                      => Sum_Nucleus_inst_mmio_bready,
      mmio_bresp                       => Sum_Nucleus_inst_mmio_bresp,
      mmio_arvalid                     => Sum_Nucleus_inst_mmio_arvalid,
      mmio_arready                     => Sum_Nucleus_inst_mmio_arready,
      mmio_araddr                      => Sum_Nucleus_inst_mmio_araddr,
      mmio_rvalid                      => Sum_Nucleus_inst_mmio_rvalid,
      mmio_rready                      => Sum_Nucleus_inst_mmio_rready,
      mmio_rdata                       => Sum_Nucleus_inst_mmio_rdata,
      mmio_rresp                       => Sum_Nucleus_inst_mmio_rresp,
      ExampleBatch_number_valid        => Sum_Nucleus_inst_ExampleBatch_number_valid,
      ExampleBatch_number_ready        => Sum_Nucleus_inst_ExampleBatch_number_ready,
      ExampleBatch_number_dvalid       => Sum_Nucleus_inst_ExampleBatch_number_dvalid,
      ExampleBatch_number_last         => Sum_Nucleus_inst_ExampleBatch_number_last,
      ExampleBatch_number              => Sum_Nucleus_inst_ExampleBatch_number,
      ExampleBatch_number_unl_valid    => Sum_Nucleus_inst_ExampleBatch_number_unl_valid,
      ExampleBatch_number_unl_ready    => Sum_Nucleus_inst_ExampleBatch_number_unl_ready,
      ExampleBatch_number_unl_tag      => Sum_Nucleus_inst_ExampleBatch_number_unl_tag,
      ExampleBatch_number_cmd_valid    => Sum_Nucleus_inst_ExampleBatch_number_cmd_valid,
      ExampleBatch_number_cmd_ready    => Sum_Nucleus_inst_ExampleBatch_number_cmd_ready,
      ExampleBatch_number_cmd_firstIdx => Sum_Nucleus_inst_ExampleBatch_number_cmd_firstIdx,
      ExampleBatch_number_cmd_lastIdx  => Sum_Nucleus_inst_ExampleBatch_number_cmd_lastIdx,
      ExampleBatch_number_cmd_ctrl     => Sum_Nucleus_inst_ExampleBatch_number_cmd_ctrl,
      ExampleBatch_number_cmd_tag      => Sum_Nucleus_inst_ExampleBatch_number_cmd_tag
    );

  Sum_ExampleBatch_inst : Sum_ExampleBatch
    generic map (
      INDEX_WIDTH                            => INDEX_WIDTH,
      TAG_WIDTH                              => TAG_WIDTH,
      EXAMPLEBATCH_NUMBER_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      EXAMPLEBATCH_NUMBER_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      EXAMPLEBATCH_NUMBER_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      EXAMPLEBATCH_NUMBER_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      EXAMPLEBATCH_NUMBER_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                            => Sum_ExampleBatch_inst_bcd_clk,
      bcd_reset                          => Sum_ExampleBatch_inst_bcd_reset,
      kcd_clk                            => Sum_ExampleBatch_inst_kcd_clk,
      kcd_reset                          => Sum_ExampleBatch_inst_kcd_reset,
      ExampleBatch_number_valid          => Sum_ExampleBatch_inst_ExampleBatch_number_valid,
      ExampleBatch_number_ready          => Sum_ExampleBatch_inst_ExampleBatch_number_ready,
      ExampleBatch_number_dvalid         => Sum_ExampleBatch_inst_ExampleBatch_number_dvalid,
      ExampleBatch_number_last           => Sum_ExampleBatch_inst_ExampleBatch_number_last,
      ExampleBatch_number                => Sum_ExampleBatch_inst_ExampleBatch_number,
      ExampleBatch_number_bus_rreq_valid => Sum_ExampleBatch_inst_ExampleBatch_number_bus_rreq_valid,
      ExampleBatch_number_bus_rreq_ready => Sum_ExampleBatch_inst_ExampleBatch_number_bus_rreq_ready,
      ExampleBatch_number_bus_rreq_addr  => Sum_ExampleBatch_inst_ExampleBatch_number_bus_rreq_addr,
      ExampleBatch_number_bus_rreq_len   => Sum_ExampleBatch_inst_ExampleBatch_number_bus_rreq_len,
      ExampleBatch_number_bus_rdat_valid => Sum_ExampleBatch_inst_ExampleBatch_number_bus_rdat_valid,
      ExampleBatch_number_bus_rdat_ready => Sum_ExampleBatch_inst_ExampleBatch_number_bus_rdat_ready,
      ExampleBatch_number_bus_rdat_data  => Sum_ExampleBatch_inst_ExampleBatch_number_bus_rdat_data,
      ExampleBatch_number_bus_rdat_last  => Sum_ExampleBatch_inst_ExampleBatch_number_bus_rdat_last,
      ExampleBatch_number_cmd_valid      => Sum_ExampleBatch_inst_ExampleBatch_number_cmd_valid,
      ExampleBatch_number_cmd_ready      => Sum_ExampleBatch_inst_ExampleBatch_number_cmd_ready,
      ExampleBatch_number_cmd_firstIdx   => Sum_ExampleBatch_inst_ExampleBatch_number_cmd_firstIdx,
      ExampleBatch_number_cmd_lastIdx    => Sum_ExampleBatch_inst_ExampleBatch_number_cmd_lastIdx,
      ExampleBatch_number_cmd_ctrl       => Sum_ExampleBatch_inst_ExampleBatch_number_cmd_ctrl,
      ExampleBatch_number_cmd_tag        => Sum_ExampleBatch_inst_ExampleBatch_number_cmd_tag,
      ExampleBatch_number_unl_valid      => Sum_ExampleBatch_inst_ExampleBatch_number_unl_valid,
      ExampleBatch_number_unl_ready      => Sum_ExampleBatch_inst_ExampleBatch_number_unl_ready,
      ExampleBatch_number_unl_tag        => Sum_ExampleBatch_inst_ExampleBatch_number_unl_tag
    );

  RDAW64DW512LW8BS1BM16_inst : BusReadArbiterVec
    generic map (
      BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH  => BUS_DATA_WIDTH,
      BUS_LEN_WIDTH   => BUS_LEN_WIDTH,
      NUM_SLAVE_PORTS => 1,
      ARB_METHOD      => "RR-STICKY",
      MAX_OUTSTANDING => 4,
      RAM_CONFIG      => "",
      SLV_REQ_SLICES  => true,
      MST_REQ_SLICE   => true,
      MST_DAT_SLICE   => true,
      SLV_DAT_SLICES  => true
    )
    port map (
      bcd_clk        => RDAW64DW512LW8BS1BM16_inst_bcd_clk,
      bcd_reset      => RDAW64DW512LW8BS1BM16_inst_bcd_reset,
      mst_rreq_valid => RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid,
      mst_rreq_ready => RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready,
      mst_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr,
      mst_rreq_len   => RDAW64DW512LW8BS1BM16_inst_mst_rreq_len,
      mst_rdat_valid => RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid,
      mst_rdat_ready => RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready,
      mst_rdat_data  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_data,
      mst_rdat_last  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_last,
      bsv_rreq_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid,
      bsv_rreq_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready,
      bsv_rreq_len   => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len,
      bsv_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr,
      bsv_rdat_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid,
      bsv_rdat_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready,
      bsv_rdat_last  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last,
      bsv_rdat_data  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data
    );

  rd_mst_rreq_valid                         <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready <= rd_mst_rreq_ready;
  rd_mst_rreq_addr                          <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr;
  rd_mst_rreq_len                           <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid <= rd_mst_rdat_valid;
  rd_mst_rdat_ready                         <= RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_data  <= rd_mst_rdat_data;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_last  <= rd_mst_rdat_last;

  Sum_Nucleus_inst_kcd_clk                               <= kcd_clk;
  Sum_Nucleus_inst_kcd_reset                             <= kcd_reset;

  Sum_Nucleus_inst_mmio_awvalid                          <= mmio_awvalid;
  mmio_awready                                           <= Sum_Nucleus_inst_mmio_awready;
  Sum_Nucleus_inst_mmio_awaddr                           <= mmio_awaddr;
  Sum_Nucleus_inst_mmio_wvalid                           <= mmio_wvalid;
  mmio_wready                                            <= Sum_Nucleus_inst_mmio_wready;
  Sum_Nucleus_inst_mmio_wdata                            <= mmio_wdata;
  Sum_Nucleus_inst_mmio_wstrb                            <= mmio_wstrb;
  mmio_bvalid                                            <= Sum_Nucleus_inst_mmio_bvalid;
  Sum_Nucleus_inst_mmio_bready                           <= mmio_bready;
  mmio_bresp                                             <= Sum_Nucleus_inst_mmio_bresp;
  Sum_Nucleus_inst_mmio_arvalid                          <= mmio_arvalid;
  mmio_arready                                           <= Sum_Nucleus_inst_mmio_arready;
  Sum_Nucleus_inst_mmio_araddr                           <= mmio_araddr;
  mmio_rvalid                                            <= Sum_Nucleus_inst_mmio_rvalid;
  Sum_Nucleus_inst_mmio_rready                           <= mmio_rready;
  mmio_rdata                                             <= Sum_Nucleus_inst_mmio_rdata;
  mmio_rresp                                             <= Sum_Nucleus_inst_mmio_rresp;

  Sum_Nucleus_inst_ExampleBatch_number_valid             <= Sum_ExampleBatch_inst_ExampleBatch_number_valid;
  Sum_ExampleBatch_inst_ExampleBatch_number_ready        <= Sum_Nucleus_inst_ExampleBatch_number_ready;
  Sum_Nucleus_inst_ExampleBatch_number_dvalid            <= Sum_ExampleBatch_inst_ExampleBatch_number_dvalid;
  Sum_Nucleus_inst_ExampleBatch_number_last              <= Sum_ExampleBatch_inst_ExampleBatch_number_last;
  Sum_Nucleus_inst_ExampleBatch_number                   <= Sum_ExampleBatch_inst_ExampleBatch_number;

  Sum_Nucleus_inst_ExampleBatch_number_unl_valid         <= Sum_ExampleBatch_inst_ExampleBatch_number_unl_valid;
  Sum_ExampleBatch_inst_ExampleBatch_number_unl_ready    <= Sum_Nucleus_inst_ExampleBatch_number_unl_ready;
  Sum_Nucleus_inst_ExampleBatch_number_unl_tag           <= Sum_ExampleBatch_inst_ExampleBatch_number_unl_tag;

  Sum_ExampleBatch_inst_bcd_clk                          <= bcd_clk;
  Sum_ExampleBatch_inst_bcd_reset                        <= bcd_reset;

  Sum_ExampleBatch_inst_kcd_clk                          <= kcd_clk;
  Sum_ExampleBatch_inst_kcd_reset                        <= kcd_reset;

  Sum_ExampleBatch_inst_ExampleBatch_number_cmd_valid    <= Sum_Nucleus_inst_ExampleBatch_number_cmd_valid;
  Sum_Nucleus_inst_ExampleBatch_number_cmd_ready         <= Sum_ExampleBatch_inst_ExampleBatch_number_cmd_ready;
  Sum_ExampleBatch_inst_ExampleBatch_number_cmd_firstIdx <= Sum_Nucleus_inst_ExampleBatch_number_cmd_firstIdx;
  Sum_ExampleBatch_inst_ExampleBatch_number_cmd_lastIdx  <= Sum_Nucleus_inst_ExampleBatch_number_cmd_lastIdx;
  Sum_ExampleBatch_inst_ExampleBatch_number_cmd_ctrl     <= Sum_Nucleus_inst_ExampleBatch_number_cmd_ctrl;
  Sum_ExampleBatch_inst_ExampleBatch_number_cmd_tag      <= Sum_Nucleus_inst_ExampleBatch_number_cmd_tag;

  RDAW64DW512LW8BS1BM16_inst_bcd_clk                     <= bcd_clk;
  RDAW64DW512LW8BS1BM16_inst_bcd_reset                   <= bcd_reset;

  Sum_ExampleBatch_inst_ExampleBatch_number_bus_rreq_ready            <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(0);
  Sum_ExampleBatch_inst_ExampleBatch_number_bus_rdat_valid            <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(0);
  Sum_ExampleBatch_inst_ExampleBatch_number_bus_rdat_last             <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(0);
  Sum_ExampleBatch_inst_ExampleBatch_number_bus_rdat_data             <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH-1 downto 0);
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(0)                        <= Sum_ExampleBatch_inst_ExampleBatch_number_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH-1 downto 0)   <= Sum_ExampleBatch_inst_ExampleBatch_number_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH-1 downto 0) <= Sum_ExampleBatch_inst_ExampleBatch_number_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(0)                        <= Sum_ExampleBatch_inst_ExampleBatch_number_bus_rdat_ready;

end architecture;
