-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Stream_pkg.all;
use work.SequenceStream_pkg.all;
use work.StreamSliceArray_pkg.all;


entity Abs_kernel is
  generic (
    INDEX_WIDTH : integer := 32;
    TAG_WIDTH   : integer := 1
  );
  port (
    kcd_clk                       : in  std_logic;
    kcd_reset                     : in  std_logic;
    BatchIn_vectors_valid         : in  std_logic;
    BatchIn_vectors_ready         : out std_logic;
    BatchIn_vectors_dvalid        : in  std_logic;
    BatchIn_vectors_last          : in  std_logic;
    BatchIn_vectors               : in  std_logic_vector(63 downto 0);
    BatchIn_vectors_unl_valid     : in  std_logic;
    BatchIn_vectors_unl_ready     : out std_logic;
    BatchIn_vectors_unl_tag       : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    BatchIn_vectors_cmd_valid     : out std_logic;
    BatchIn_vectors_cmd_ready     : in  std_logic;
    BatchIn_vectors_cmd_firstIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    BatchIn_vectors_cmd_lastIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    BatchIn_vectors_cmd_tag       : out std_logic_vector(TAG_WIDTH-1 downto 0);
    BatchOut_vectors_valid        : out std_logic;
    BatchOut_vectors_ready        : in  std_logic;
    BatchOut_vectors_dvalid       : out std_logic := '1';
    BatchOut_vectors_last         : out std_logic;
    BatchOut_vectors              : out std_logic_vector(63 downto 0);
    BatchOut_vectors_unl_valid    : in  std_logic;
    BatchOut_vectors_unl_ready    : out std_logic;
    BatchOut_vectors_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    BatchOut_vectors_cmd_valid    : out std_logic;
    BatchOut_vectors_cmd_ready    : in  std_logic;
    BatchOut_vectors_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    BatchOut_vectors_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    BatchOut_vectors_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    start                         : in  std_logic;
    stop                          : in  std_logic;
    reset                         : in  std_logic;
    idle                          : out std_logic;
    busy                          : out std_logic;
    done                          : out std_logic;
    result                        : out std_logic_vector(63 downto 0);
    BatchIn_firstidx              : in  std_logic_vector(31 downto 0);
    BatchIn_lastidx               : in  std_logic_vector(31 downto 0);
    BatchOut_firstidx             : in  std_logic_vector(31 downto 0);
    BatchOut_lastidx              : in  std_logic_vector(31 downto 0)
  );
end entity;

architecture Implementation of Abs_kernel is

  signal count_valid                : std_logic;
  signal count_ready                : std_logic;
  signal count                      : std_logic_vector(8-1 downto 0);
  signal count_last                 : std_logic;
  
  
  
  signal counter_valid              : std_logic;
  signal counter_ready              : std_logic;
  
  signal seq_valid                  : std_logic;
  signal seq_ready                  : std_logic;
  
  signal dly_in_valid               :std_logic;
  signal dly_in_ready               :std_logic;
  signal dly_in_data                : std_logic_vector(63 downto 0);
  
  signal dly_out_valid               :std_logic;
  signal dly_out_ready               :std_logic;
  signal dly_out_data                :std_logic_vector(63 downto 0);
  
  
  -- Enumeration type for our state machine.
  type state_t is (STATE_IDLE, 
                   STATE_COMMAND, 
                   STATE_CALCULATING, 
                   STATE_UNLOCK, 
                   STATE_DONE);
  
  -- Current state register and next state signal.
	signal state, state_next : state_t;

begin

element_counter: StreamElementCounter
    generic map (
      IN_COUNT_MAX              => 10,
      IN_COUNT_WIDTH            => 8,
      OUT_COUNT_MAX             => 10,
      OUT_COUNT_WIDTH           => 8
    )
    port map (
      clk                       => kcd_clk,
      reset                     => reset,
      in_valid                  => counter_valid,
      in_ready                  => counter_ready,
      in_dvalid                 => BatchIn_vectors_dvalid,
      in_count                  => "00000001",
      in_last                   => BatchIn_vectors_last,
      out_valid                 => count_valid,
      out_ready                 => count_ready,
      out_last                  => count_last,
      out_count                 => count
    );
    
    
 sequencer: SequenceStream
    generic map (
      MIN_BUFFER_DEPTH           => 10,
      LENGTH_WIDTH               => 8,
      BLOCKING                   => false
    )
    port map (
      clk                       => kcd_clk,
      reset                     => reset,
      in_valid                  => dly_out_valid,
      in_ready                  => dly_out_ready,
      in_dvalid                 => '1',
      in_count                  => "00000001",
      in_length_valid           => count_valid,
      in_length_ready           => count_ready,
      in_length_data            => count,
      out_valid                 => BatchOut_vectors_valid,
      out_ready                 => BatchOut_vectors_ready,
      out_last                  => BatchOut_vectors_last
    );
    
    --Connect data lanes outside the module
    
    BatchOut_vectors <= dly_out_data;
    
    dly: StreamSliceArray
    generic map (
      DATA_WIDTH                 => 64,
      DEPTH                      => 10
    )
    port map (
      clk                       => kcd_clk,
      reset                     => reset,

      in_valid                  => dly_in_valid,
      in_ready                  => dly_in_ready,
      in_data                   => BatchIn_vectors,

      out_valid                 => dly_out_valid,
      out_ready                 => dly_out_ready,
      out_data                  => dly_out_data

    );
    
    sync: StreamSync
    generic map (
      NUM_INPUTS                => 1,
      NUM_OUTPUTS               => 2
    )
    port map (
      clk                       => kcd_clk,
      reset                     => reset,

      in_valid(0)               => BatchIn_vectors_valid,
      in_ready(0)               => BatchIn_vectors_ready,


      out_valid(0)              => counter_valid,
      out_valid(1)              => dly_in_valid,
      out_ready(0)              => counter_ready,
      out_ready(1)              => dly_in_ready

    );

    

  combinatorial_proc : process (all) is 
  begin
    
    -- We first determine the default outputs of our combinatorial circuit.
    -- They may be overwritten by sequential statements within this process
    -- later on.
    
    -- Make sure the command stream is deasserted by default.
    BatchIn_vectors_cmd_valid    <= '0';
    BatchIn_vectors_cmd_firstIdx <= (others => '0');
    BatchIn_vectors_cmd_lastIdx  <= (others => '0');
    BatchIn_vectors_cmd_tag      <= (others => '0');
    
    BatchOut_vectors_cmd_valid    <= '0';
    BatchOut_vectors_cmd_firstIdx <= (others => '0');
    BatchOut_vectors_cmd_lastIdx  <= (others => '0');
    BatchOut_vectors_cmd_tag      <= (others => '0');
    
    BatchIn_vectors_unl_ready <= '0'; -- Do not accept "unlocks".
    state_next <= state;                  -- Retain current state.

    -- For every state, we will determine the outputs of our combinatorial 
    -- circuit.
    case state is
      when STATE_IDLE =>
        -- Idle: We just wait for the start bit to come up.
        done <= '0';
        busy <= '0';
        idle <= '1';
                
        -- Wait for the start signal (typically controlled by the host-side 
        -- software).
        if start = '1' then
          state_next <= STATE_COMMAND;
        end if;

      when STATE_COMMAND =>
        -- Command: we send a command to the generated interface.
        done <= '0';
        busy <= '1';  
        idle <= '0';
                
        -- The command is a stream, so we assert its valid bit and wait in this
        -- state until it is accepted by the generated interface. If the valid
        -- and ready bit are both asserted in the same cycle, the command is
        -- accepted.        
        -- We need to supply a command to the generated interface for each 
        -- Arrow field. In the case of this kernel, that means we just have to
        -- generate a single command. The command is sent on the command stream 
        -- to the generated interface.
        -- The command includes a range of rows from the recordbatch we want to
        -- work on. In this simple example, we just want this kernel to work on 
        -- all the rows in the RecordBatch. 
        -- The starting row and ending row (exclusive) that this kernel should 
        -- work on is supplied via MMIO and appears on the firstIdx and lastIdx 
        -- ports.
        -- We can use the tag field of the command stream to identify different 
        -- commands. We don't really use it for this example, so we just set it
        -- to zero.
        BatchIn_vectors_cmd_valid    <= '1';
        BatchIn_vectors_cmd_firstIdx <= BatchIn_firstIdx;
        BatchIn_vectors_cmd_lastIdx  <= BatchIn_lastIdx;
        BatchIn_vectors_cmd_tag      <= (others => '0');
        
        Batchout_vectors_cmd_valid    <= '1';
        BatchOut_vectors_cmd_firstIdx <= BatchIn_firstIdx;
        BatchOut_vectors_cmd_lastIdx  <= BatchIn_lastIdx;
        BatchOut_vectors_cmd_tag      <= (others => '0');
        
        if BatchIn_vectors_cmd_ready = '1' and BatchOut_vectors_cmd_ready = '1' then
          state_next <= STATE_CALCULATING;
        end if;

      when STATE_CALCULATING =>
        -- Calculating: we stream in and accumulate the numbers one by one.
        done <= '0';
        busy <= '1';  
        idle <= '0';
          
          -- All we have to do now is check if the last number was supplied.
          -- If that is the case, we can go to the "done" state.
          if BatchOut_vectors_last = '1' then
            state_next <= STATE_UNLOCK;
          end if;
        
      when STATE_UNLOCK =>
        -- Unlock: the generated interface delivered all items in the stream.
        -- The unlock stream is supplied to make sure all bus transfers of the
        -- corresponding command are completed.
        done <= '1';
        busy <= '0';
        idle <= '1';
        
        -- Ready to handshake the unlock stream:
        BatchIn_vectors_unl_ready <= '1';
        Batchout_vectors_unl_ready <= '1';
        -- Handshake when it is valid and go to the done state.
        if BatchIn_vectors_unl_valid = '1' and BatchOut_vectors_unl_valid = '1' then
          state_next <= STATE_DONE;
        end if;

      when STATE_DONE =>
        -- Done: the kernel is done with its job.
        done <= '1';
        busy <= '0';
        idle <= '1';
        
        -- Wait for the reset signal (typically controlled by the host-side 
        -- software), so we can go to idle again. This reset is not to be
        -- confused with the system-wide reset that travels into the kernel
        -- alongside the clock (kcd_reset).
        if reset = '1' then
          state_next <= STATE_IDLE;
        end if;
        
    end case;
  end process;


 -- Sequential part:
  sequential_proc: process (kcd_clk)
  begin
    -- On the rising edge of the kernel clock:
    if rising_edge(kcd_clk) then
      -- Register the next state.
      state <= state_next;
        
      -- If there is a (synchronous) reset, go to idle and make the 
      -- accumulator hold zero.
      if kcd_reset = '1' then
        state <= STATE_IDLE;
      end if;
    end if;
  end process;

end architecture;
