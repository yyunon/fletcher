-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;

entity Abs_kernel_BatchOut is
  generic (
    INDEX_WIDTH                         : integer := 32;
    TAG_WIDTH                           : integer := 1;
    BATCHOUT_VECTORS_BUS_ADDR_WIDTH     : integer := 64;
    BATCHOUT_VECTORS_BUS_DATA_WIDTH     : integer := 512;
    BATCHOUT_VECTORS_BUS_LEN_WIDTH      : integer := 8;
    BATCHOUT_VECTORS_BUS_BURST_STEP_LEN : integer := 1;
    BATCHOUT_VECTORS_BUS_BURST_MAX_LEN  : integer := 16
  );
  port (
    bcd_clk                          : in  std_logic;
    bcd_reset                        : in  std_logic;
    kcd_clk                          : in  std_logic;
    kcd_reset                        : in  std_logic;
    BatchOut_vectors_valid           : in  std_logic;
    BatchOut_vectors_ready           : out std_logic;
    BatchOut_vectors_dvalid          : in  std_logic;
    BatchOut_vectors_last            : in  std_logic;
    BatchOut_vectors                 : in  std_logic_vector(63 downto 0);
    BatchOut_vectors_bus_wreq_valid  : out std_logic;
    BatchOut_vectors_bus_wreq_ready  : in  std_logic;
    BatchOut_vectors_bus_wreq_addr   : out std_logic_vector(BATCHOUT_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
    BatchOut_vectors_bus_wreq_len    : out std_logic_vector(BATCHOUT_VECTORS_BUS_LEN_WIDTH-1 downto 0);
    BatchOut_vectors_bus_wdat_valid  : out std_logic;
    BatchOut_vectors_bus_wdat_ready  : in  std_logic;
    BatchOut_vectors_bus_wdat_data   : out std_logic_vector(BATCHOUT_VECTORS_BUS_DATA_WIDTH-1 downto 0);
    BatchOut_vectors_bus_wdat_strobe : out std_logic_vector(BATCHOUT_VECTORS_BUS_DATA_WIDTH/8-1 downto 0);
    BatchOut_vectors_bus_wdat_last   : out std_logic;
    BatchOut_vectors_cmd_valid       : in  std_logic;
    BatchOut_vectors_cmd_ready       : out std_logic;
    BatchOut_vectors_cmd_firstIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    BatchOut_vectors_cmd_lastIdx     : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    BatchOut_vectors_cmd_ctrl        : in  std_logic_vector(BATCHOUT_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
    BatchOut_vectors_cmd_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    BatchOut_vectors_unl_valid       : out std_logic;
    BatchOut_vectors_unl_ready       : in  std_logic;
    BatchOut_vectors_unl_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0)
  );
end entity;

architecture Implementation of Abs_kernel_BatchOut is
  signal vectors_inst_bcd_clk         : std_logic;
  signal vectors_inst_bcd_reset       : std_logic;

  signal vectors_inst_kcd_clk         : std_logic;
  signal vectors_inst_kcd_reset       : std_logic;

  signal vectors_inst_cmd_valid       : std_logic;
  signal vectors_inst_cmd_ready       : std_logic;
  signal vectors_inst_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal vectors_inst_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal vectors_inst_cmd_ctrl        : std_logic_vector(BATCHOUT_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
  signal vectors_inst_cmd_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal vectors_inst_unl_valid       : std_logic;
  signal vectors_inst_unl_ready       : std_logic;
  signal vectors_inst_unl_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal vectors_inst_bus_wreq_valid  : std_logic;
  signal vectors_inst_bus_wreq_ready  : std_logic;
  signal vectors_inst_bus_wreq_addr   : std_logic_vector(BATCHOUT_VECTORS_BUS_ADDR_WIDTH-1 downto 0);
  signal vectors_inst_bus_wreq_len    : std_logic_vector(BATCHOUT_VECTORS_BUS_LEN_WIDTH-1 downto 0);
  signal vectors_inst_bus_wdat_valid  : std_logic;
  signal vectors_inst_bus_wdat_ready  : std_logic;
  signal vectors_inst_bus_wdat_data   : std_logic_vector(BATCHOUT_VECTORS_BUS_DATA_WIDTH-1 downto 0);
  signal vectors_inst_bus_wdat_strobe : std_logic_vector(BATCHOUT_VECTORS_BUS_DATA_WIDTH/8-1 downto 0);
  signal vectors_inst_bus_wdat_last   : std_logic;

  signal vectors_inst_in_valid        : std_logic_vector(0 downto 0);
  signal vectors_inst_in_ready        : std_logic_vector(0 downto 0);
  signal vectors_inst_in_data         : std_logic_vector(63 downto 0);
  signal vectors_inst_in_dvalid       : std_logic_vector(0 downto 0);
  signal vectors_inst_in_last         : std_logic_vector(0 downto 0);

begin
  vectors_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH     => BATCHOUT_VECTORS_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => BATCHOUT_VECTORS_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => BATCHOUT_VECTORS_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => BATCHOUT_VECTORS_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => BATCHOUT_VECTORS_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk         => vectors_inst_bcd_clk,
      bcd_reset       => vectors_inst_bcd_reset,
      kcd_clk         => vectors_inst_kcd_clk,
      kcd_reset       => vectors_inst_kcd_reset,
      cmd_valid       => vectors_inst_cmd_valid,
      cmd_ready       => vectors_inst_cmd_ready,
      cmd_firstIdx    => vectors_inst_cmd_firstIdx,
      cmd_lastIdx     => vectors_inst_cmd_lastIdx,
      cmd_ctrl        => vectors_inst_cmd_ctrl,
      cmd_tag         => vectors_inst_cmd_tag,
      unl_valid       => vectors_inst_unl_valid,
      unl_ready       => vectors_inst_unl_ready,
      unl_tag         => vectors_inst_unl_tag,
      bus_wreq_valid  => vectors_inst_bus_wreq_valid,
      bus_wreq_ready  => vectors_inst_bus_wreq_ready,
      bus_wreq_addr   => vectors_inst_bus_wreq_addr,
      bus_wreq_len    => vectors_inst_bus_wreq_len,
      bus_wdat_valid  => vectors_inst_bus_wdat_valid,
      bus_wdat_ready  => vectors_inst_bus_wdat_ready,
      bus_wdat_data   => vectors_inst_bus_wdat_data,
      bus_wdat_strobe => vectors_inst_bus_wdat_strobe,
      bus_wdat_last   => vectors_inst_bus_wdat_last,
      in_valid        => vectors_inst_in_valid,
      in_ready        => vectors_inst_in_ready,
      in_data         => vectors_inst_in_data,
      in_dvalid       => vectors_inst_in_dvalid,
      in_last         => vectors_inst_in_last
    );

  BatchOut_vectors_bus_wreq_valid  <= vectors_inst_bus_wreq_valid;
  vectors_inst_bus_wreq_ready      <= BatchOut_vectors_bus_wreq_ready;
  BatchOut_vectors_bus_wreq_addr   <= vectors_inst_bus_wreq_addr;
  BatchOut_vectors_bus_wreq_len    <= vectors_inst_bus_wreq_len;
  BatchOut_vectors_bus_wdat_valid  <= vectors_inst_bus_wdat_valid;
  vectors_inst_bus_wdat_ready      <= BatchOut_vectors_bus_wdat_ready;
  BatchOut_vectors_bus_wdat_data   <= vectors_inst_bus_wdat_data;
  BatchOut_vectors_bus_wdat_strobe <= vectors_inst_bus_wdat_strobe;
  BatchOut_vectors_bus_wdat_last   <= vectors_inst_bus_wdat_last;

  BatchOut_vectors_unl_valid       <= vectors_inst_unl_valid;
  vectors_inst_unl_ready           <= BatchOut_vectors_unl_ready;
  BatchOut_vectors_unl_tag         <= vectors_inst_unl_tag;

  vectors_inst_bcd_clk       <= bcd_clk;
  vectors_inst_bcd_reset     <= bcd_reset;

  vectors_inst_kcd_clk       <= kcd_clk;
  vectors_inst_kcd_reset     <= kcd_reset;

  vectors_inst_cmd_valid     <= BatchOut_vectors_cmd_valid;
  BatchOut_vectors_cmd_ready <= vectors_inst_cmd_ready;
  vectors_inst_cmd_firstIdx  <= BatchOut_vectors_cmd_firstIdx;
  vectors_inst_cmd_lastIdx   <= BatchOut_vectors_cmd_lastIdx;
  vectors_inst_cmd_ctrl      <= BatchOut_vectors_cmd_ctrl;
  vectors_inst_cmd_tag       <= BatchOut_vectors_cmd_tag;

  vectors_inst_in_valid(0)   <= BatchOut_vectors_valid;
  BatchOut_vectors_ready     <= vectors_inst_in_ready(0);
  vectors_inst_in_data       <= BatchOut_vectors;
  vectors_inst_in_dvalid(0)  <= BatchOut_vectors_dvalid;
  vectors_inst_in_last(0)    <= BatchOut_vectors_last;

end architecture;
