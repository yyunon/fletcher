-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;
use work.mmio_pkg.all;

entity Sum_Nucleus is
  generic (
    INDEX_WIDTH                        : integer := 32;
    TAG_WIDTH                          : integer := 1;
    EXAMPLEBATCH_NUMBER_BUS_ADDR_WIDTH : integer := 64
  );
  port (
    kcd_clk                          : in  std_logic;
    kcd_reset                        : in  std_logic;
    mmio_awvalid                     : in  std_logic;
    mmio_awready                     : out std_logic;
    mmio_awaddr                      : in  std_logic_vector(31 downto 0);
    mmio_wvalid                      : in  std_logic;
    mmio_wready                      : out std_logic;
    mmio_wdata                       : in  std_logic_vector(31 downto 0);
    mmio_wstrb                       : in  std_logic_vector(3 downto 0);
    mmio_bvalid                      : out std_logic;
    mmio_bready                      : in  std_logic;
    mmio_bresp                       : out std_logic_vector(1 downto 0);
    mmio_arvalid                     : in  std_logic;
    mmio_arready                     : out std_logic;
    mmio_araddr                      : in  std_logic_vector(31 downto 0);
    mmio_rvalid                      : out std_logic;
    mmio_rready                      : in  std_logic;
    mmio_rdata                       : out std_logic_vector(31 downto 0);
    mmio_rresp                       : out std_logic_vector(1 downto 0);
    ExampleBatch_number_valid        : in  std_logic;
    ExampleBatch_number_ready        : out std_logic;
    ExampleBatch_number_dvalid       : in  std_logic;
    ExampleBatch_number_last         : in  std_logic;
    ExampleBatch_number              : in  std_logic_vector(63 downto 0);
    ExampleBatch_number_unl_valid    : in  std_logic;
    ExampleBatch_number_unl_ready    : out std_logic;
    ExampleBatch_number_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ExampleBatch_number_cmd_valid    : out std_logic;
    ExampleBatch_number_cmd_ready    : in  std_logic;
    ExampleBatch_number_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ExampleBatch_number_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ExampleBatch_number_cmd_ctrl     : out std_logic_vector(EXAMPLEBATCH_NUMBER_BUS_ADDR_WIDTH-1 downto 0);
    ExampleBatch_number_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0)
  );
end entity;

architecture Implementation of Sum_Nucleus is
  component Sum is
    generic (
      INDEX_WIDTH : integer := 32;
      TAG_WIDTH   : integer := 1
    );
    port (
      kcd_clk                          : in  std_logic;
      kcd_reset                        : in  std_logic;
      ExampleBatch_number_valid        : in  std_logic;
      ExampleBatch_number_ready        : out std_logic;
      ExampleBatch_number_dvalid       : in  std_logic;
      ExampleBatch_number_last         : in  std_logic;
      ExampleBatch_number              : in  std_logic_vector(63 downto 0);
      ExampleBatch_number_unl_valid    : in  std_logic;
      ExampleBatch_number_unl_ready    : out std_logic;
      ExampleBatch_number_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ExampleBatch_number_cmd_valid    : out std_logic;
      ExampleBatch_number_cmd_ready    : in  std_logic;
      ExampleBatch_number_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ExampleBatch_number_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ExampleBatch_number_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      start                            : in  std_logic;
      stop                             : in  std_logic;
      reset                            : in  std_logic;
      idle                             : out std_logic;
      busy                             : out std_logic;
      done                             : out std_logic;
      result                           : out std_logic_vector(63 downto 0);
      ExampleBatch_firstidx            : in  std_logic_vector(31 downto 0);
      ExampleBatch_lastidx             : in  std_logic_vector(31 downto 0)
    );
  end component;

  signal Sum_inst_kcd_clk                                       : std_logic;
  signal Sum_inst_kcd_reset                                     : std_logic;

  signal Sum_inst_ExampleBatch_number_valid                     : std_logic;
  signal Sum_inst_ExampleBatch_number_ready                     : std_logic;
  signal Sum_inst_ExampleBatch_number_dvalid                    : std_logic;
  signal Sum_inst_ExampleBatch_number_last                      : std_logic;
  signal Sum_inst_ExampleBatch_number                           : std_logic_vector(63 downto 0);

  signal Sum_inst_ExampleBatch_number_unl_valid                 : std_logic;
  signal Sum_inst_ExampleBatch_number_unl_ready                 : std_logic;
  signal Sum_inst_ExampleBatch_number_unl_tag                   : std_logic_vector(0 downto 0);

  signal Sum_inst_ExampleBatch_number_cmd_valid                 : std_logic;
  signal Sum_inst_ExampleBatch_number_cmd_ready                 : std_logic;
  signal Sum_inst_ExampleBatch_number_cmd_firstIdx              : std_logic_vector(31 downto 0);
  signal Sum_inst_ExampleBatch_number_cmd_lastIdx               : std_logic_vector(31 downto 0);
  signal Sum_inst_ExampleBatch_number_cmd_tag                   : std_logic_vector(0 downto 0);

  signal Sum_inst_start                                         : std_logic;
  signal Sum_inst_stop                                          : std_logic;
  signal Sum_inst_reset                                         : std_logic;
  signal Sum_inst_idle                                          : std_logic;
  signal Sum_inst_busy                                          : std_logic;
  signal Sum_inst_done                                          : std_logic;
  signal Sum_inst_result                                        : std_logic_vector(63 downto 0);
  signal Sum_inst_ExampleBatch_firstidx                         : std_logic_vector(31 downto 0);
  signal Sum_inst_ExampleBatch_lastidx                          : std_logic_vector(31 downto 0);
  signal mmio_inst_kcd_clk                                      : std_logic;
  signal mmio_inst_kcd_reset                                    : std_logic;

  signal mmio_inst_f_start_data                                 : std_logic;
  signal mmio_inst_f_stop_data                                  : std_logic;
  signal mmio_inst_f_reset_data                                 : std_logic;
  signal mmio_inst_f_idle_write_data                            : std_logic;
  signal mmio_inst_f_busy_write_data                            : std_logic;
  signal mmio_inst_f_done_write_data                            : std_logic;
  signal mmio_inst_f_result_write_data                          : std_logic_vector(63 downto 0);
  signal mmio_inst_f_ExampleBatch_firstidx_data                 : std_logic_vector(31 downto 0);
  signal mmio_inst_f_ExampleBatch_lastidx_data                  : std_logic_vector(31 downto 0);
  signal mmio_inst_f_ExampleBatch_number_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_Profile_enable_data                        : std_logic;
  signal mmio_inst_f_Profile_clear_data                         : std_logic;
  signal mmio_inst_mmio_awvalid                                 : std_logic;
  signal mmio_inst_mmio_awready                                 : std_logic;
  signal mmio_inst_mmio_awaddr                                  : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wvalid                                  : std_logic;
  signal mmio_inst_mmio_wready                                  : std_logic;
  signal mmio_inst_mmio_wdata                                   : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wstrb                                   : std_logic_vector(3 downto 0);
  signal mmio_inst_mmio_bvalid                                  : std_logic;
  signal mmio_inst_mmio_bready                                  : std_logic;
  signal mmio_inst_mmio_bresp                                   : std_logic_vector(1 downto 0);
  signal mmio_inst_mmio_arvalid                                 : std_logic;
  signal mmio_inst_mmio_arready                                 : std_logic;
  signal mmio_inst_mmio_araddr                                  : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rvalid                                  : std_logic;
  signal mmio_inst_mmio_rready                                  : std_logic;
  signal mmio_inst_mmio_rdata                                   : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rresp                                   : std_logic_vector(1 downto 0);

  signal ExampleBatch_number_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal ExampleBatch_number_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal ExampleBatch_number_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ExampleBatch_number_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ExampleBatch_number_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ExampleBatch_number_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal ExampleBatch_number_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal ExampleBatch_number_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ExampleBatch_number_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ExampleBatch_number_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(EXAMPLEBATCH_NUMBER_BUS_ADDR_WIDTH-1 downto 0);
  signal ExampleBatch_number_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ExampleBatch_number_cmd_accm_inst_ctrl : std_logic_vector(EXAMPLEBATCH_NUMBER_BUS_ADDR_WIDTH-1 downto 0);

begin
  Sum_inst : Sum
    generic map (
      INDEX_WIDTH => 32,
      TAG_WIDTH   => 1
    )
    port map (
      kcd_clk                          => Sum_inst_kcd_clk,
      kcd_reset                        => Sum_inst_kcd_reset,
      ExampleBatch_number_valid        => Sum_inst_ExampleBatch_number_valid,
      ExampleBatch_number_ready        => Sum_inst_ExampleBatch_number_ready,
      ExampleBatch_number_dvalid       => Sum_inst_ExampleBatch_number_dvalid,
      ExampleBatch_number_last         => Sum_inst_ExampleBatch_number_last,
      ExampleBatch_number              => Sum_inst_ExampleBatch_number,
      ExampleBatch_number_unl_valid    => Sum_inst_ExampleBatch_number_unl_valid,
      ExampleBatch_number_unl_ready    => Sum_inst_ExampleBatch_number_unl_ready,
      ExampleBatch_number_unl_tag      => Sum_inst_ExampleBatch_number_unl_tag,
      ExampleBatch_number_cmd_valid    => Sum_inst_ExampleBatch_number_cmd_valid,
      ExampleBatch_number_cmd_ready    => Sum_inst_ExampleBatch_number_cmd_ready,
      ExampleBatch_number_cmd_firstIdx => Sum_inst_ExampleBatch_number_cmd_firstIdx,
      ExampleBatch_number_cmd_lastIdx  => Sum_inst_ExampleBatch_number_cmd_lastIdx,
      ExampleBatch_number_cmd_tag      => Sum_inst_ExampleBatch_number_cmd_tag,
      start                            => Sum_inst_start,
      stop                             => Sum_inst_stop,
      reset                            => Sum_inst_reset,
      idle                             => Sum_inst_idle,
      busy                             => Sum_inst_busy,
      done                             => Sum_inst_done,
      result                           => Sum_inst_result,
      ExampleBatch_firstidx            => Sum_inst_ExampleBatch_firstidx,
      ExampleBatch_lastidx             => Sum_inst_ExampleBatch_lastidx
    );

  mmio_inst : mmio
    port map (
      kcd_clk                           => mmio_inst_kcd_clk,
      kcd_reset                         => mmio_inst_kcd_reset,
      f_start_data                      => mmio_inst_f_start_data,
      f_stop_data                       => mmio_inst_f_stop_data,
      f_reset_data                      => mmio_inst_f_reset_data,
      f_idle_write_data                 => mmio_inst_f_idle_write_data,
      f_busy_write_data                 => mmio_inst_f_busy_write_data,
      f_done_write_data                 => mmio_inst_f_done_write_data,
      f_result_write_data               => mmio_inst_f_result_write_data,
      f_ExampleBatch_firstidx_data      => mmio_inst_f_ExampleBatch_firstidx_data,
      f_ExampleBatch_lastidx_data       => mmio_inst_f_ExampleBatch_lastidx_data,
      f_ExampleBatch_number_values_data => mmio_inst_f_ExampleBatch_number_values_data,
      mmio_awvalid                      => mmio_inst_mmio_awvalid,
      mmio_awready                      => mmio_inst_mmio_awready,
      mmio_awaddr                       => mmio_inst_mmio_awaddr,
      mmio_wvalid                       => mmio_inst_mmio_wvalid,
      mmio_wready                       => mmio_inst_mmio_wready,
      mmio_wdata                        => mmio_inst_mmio_wdata,
      mmio_wstrb                        => mmio_inst_mmio_wstrb,
      mmio_bvalid                       => mmio_inst_mmio_bvalid,
      mmio_bready                       => mmio_inst_mmio_bready,
      mmio_bresp                        => mmio_inst_mmio_bresp,
      mmio_arvalid                      => mmio_inst_mmio_arvalid,
      mmio_arready                      => mmio_inst_mmio_arready,
      mmio_araddr                       => mmio_inst_mmio_araddr,
      mmio_rvalid                       => mmio_inst_mmio_rvalid,
      mmio_rready                       => mmio_inst_mmio_rready,
      mmio_rdata                        => mmio_inst_mmio_rdata,
      mmio_rresp                        => mmio_inst_mmio_rresp
    );

  ExampleBatch_number_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => EXAMPLEBATCH_NUMBER_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => ExampleBatch_number_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => ExampleBatch_number_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => ExampleBatch_number_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => ExampleBatch_number_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => ExampleBatch_number_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => ExampleBatch_number_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => ExampleBatch_number_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => ExampleBatch_number_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => ExampleBatch_number_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => ExampleBatch_number_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => ExampleBatch_number_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => ExampleBatch_number_cmd_accm_inst_ctrl
    );

  ExampleBatch_number_cmd_valid                       <= ExampleBatch_number_cmd_accm_inst_nucleus_cmd_valid;
  ExampleBatch_number_cmd_accm_inst_nucleus_cmd_ready <= ExampleBatch_number_cmd_ready;
  ExampleBatch_number_cmd_firstIdx                    <= ExampleBatch_number_cmd_accm_inst_nucleus_cmd_firstIdx;
  ExampleBatch_number_cmd_lastIdx                     <= ExampleBatch_number_cmd_accm_inst_nucleus_cmd_lastIdx;
  ExampleBatch_number_cmd_ctrl                        <= ExampleBatch_number_cmd_accm_inst_nucleus_cmd_ctrl;
  ExampleBatch_number_cmd_tag                         <= ExampleBatch_number_cmd_accm_inst_nucleus_cmd_tag;

  Sum_inst_kcd_clk                                      <= kcd_clk;
  Sum_inst_kcd_reset                                    <= kcd_reset;

  Sum_inst_ExampleBatch_number_valid                    <= ExampleBatch_number_valid;
  ExampleBatch_number_ready                             <= Sum_inst_ExampleBatch_number_ready;
  Sum_inst_ExampleBatch_number_dvalid                   <= ExampleBatch_number_dvalid;
  Sum_inst_ExampleBatch_number_last                     <= ExampleBatch_number_last;
  Sum_inst_ExampleBatch_number                          <= ExampleBatch_number;

  Sum_inst_ExampleBatch_number_unl_valid                <= ExampleBatch_number_unl_valid;
  ExampleBatch_number_unl_ready                         <= Sum_inst_ExampleBatch_number_unl_ready;
  Sum_inst_ExampleBatch_number_unl_tag                  <= ExampleBatch_number_unl_tag;

  Sum_inst_start                                        <= mmio_inst_f_start_data;
  Sum_inst_stop                                         <= mmio_inst_f_stop_data;
  Sum_inst_reset                                        <= mmio_inst_f_reset_data;
  Sum_inst_ExampleBatch_firstidx                        <= mmio_inst_f_ExampleBatch_firstidx_data;
  Sum_inst_ExampleBatch_lastidx                         <= mmio_inst_f_ExampleBatch_lastidx_data;
  mmio_inst_kcd_clk                                     <= kcd_clk;
  mmio_inst_kcd_reset                                   <= kcd_reset;

  mmio_inst_f_idle_write_data                           <= Sum_inst_idle;
  mmio_inst_f_busy_write_data                           <= Sum_inst_busy;
  mmio_inst_f_done_write_data                           <= Sum_inst_done;
  mmio_inst_f_result_write_data                         <= Sum_inst_result;
  mmio_inst_mmio_awvalid                                <= mmio_awvalid;
  mmio_awready                                          <= mmio_inst_mmio_awready;
  mmio_inst_mmio_awaddr                                 <= mmio_awaddr;
  mmio_inst_mmio_wvalid                                 <= mmio_wvalid;
  mmio_wready                                           <= mmio_inst_mmio_wready;
  mmio_inst_mmio_wdata                                  <= mmio_wdata;
  mmio_inst_mmio_wstrb                                  <= mmio_wstrb;
  mmio_bvalid                                           <= mmio_inst_mmio_bvalid;
  mmio_inst_mmio_bready                                 <= mmio_bready;
  mmio_bresp                                            <= mmio_inst_mmio_bresp;
  mmio_inst_mmio_arvalid                                <= mmio_arvalid;
  mmio_arready                                          <= mmio_inst_mmio_arready;
  mmio_inst_mmio_araddr                                 <= mmio_araddr;
  mmio_rvalid                                           <= mmio_inst_mmio_rvalid;
  mmio_inst_mmio_rready                                 <= mmio_rready;
  mmio_rdata                                            <= mmio_inst_mmio_rdata;
  mmio_rresp                                            <= mmio_inst_mmio_rresp;

  ExampleBatch_number_cmd_accm_inst_kernel_cmd_valid    <= Sum_inst_ExampleBatch_number_cmd_valid;
  Sum_inst_ExampleBatch_number_cmd_ready                <= ExampleBatch_number_cmd_accm_inst_kernel_cmd_ready;
  ExampleBatch_number_cmd_accm_inst_kernel_cmd_firstIdx <= Sum_inst_ExampleBatch_number_cmd_firstIdx;
  ExampleBatch_number_cmd_accm_inst_kernel_cmd_lastIdx  <= Sum_inst_ExampleBatch_number_cmd_lastIdx;
  ExampleBatch_number_cmd_accm_inst_kernel_cmd_tag      <= Sum_inst_ExampleBatch_number_cmd_tag;

  ExampleBatch_number_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_ExampleBatch_number_values_data;

end architecture;
